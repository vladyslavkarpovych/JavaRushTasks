���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.5.1�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK*�verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak��ST_Slope�et�b�n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJf��_hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��h3�f8�����R�(KhQNNNJ����J����K t�b�C              �?�t�bhUh'�scalar���hPC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hK�
node_count�Kٌnodes�h)h,K ��h.��R�(KKم�h3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h�hPK ��h�hPK��h�hPK��h�hbK��h�hbK ��h�hPK(��h�hbK0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@6         ^       	          033�?���:���?�           ��@                                 �_@z�t���?�             x@                                   �?D|U��@�?.            �P@                                  �?���?            �D@                                 �_@���Q��?             9@              	                   �[@�t����?	             1@                                  �`@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        
                          `]@ףp=
�?             $@        ������������������������       �                     @                      
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   @K@      �?              @                                  �\@      �?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �                     :@               C                    �?l�"���?�            �s@               :                    �?��7	C)�?D            @Z@              !                     D@���o,��?.            @R@                                   �B@      �?              @        ������������������������       �                     �?                                   Hq@؇���X�?             @                                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        "       '                   �_@؇>���?)            @P@        #       &       
             �?�\��N��?             3@       $       %                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     "@        (       -                    �?*
;&���?             G@        )       ,                    b@���|���?             &@       *       +                   `\@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        .       /                   �l@�#-���?            �A@        ������������������������       �        
             5@        0       1                   �Z@d}h���?             ,@        ������������������������       �                     �?        2       9       	          ����?8�Z$���?
             *@       3       4                   �m@"pc�
�?             &@        ������������������������       �                     �?        5       6                   �a@ףp=
�?             $@       ������������������������       �                     @        7       8                    d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ;       >       
             �?     ��?             @@       <       =                   �b@ףp=
�?             4@       ������������������������       �                     2@        ������������������������       �                      @        ?       @                   �a@�q�q�?             (@        ������������������������       �                     @        A       B                   �^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        D       S       
             �?@mW���?�            �j@        E       J                    �J@�K��&�?            �E@        F       G                    �?�<ݚ�?             2@       ������������������������       �                     *@        H       I                    @E@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        K       L                    �?�J�4�?             9@        ������������������������       �                     �?        M       R                   �l@      �?             8@        N       O                    �?      �?              @        ������������������������       �                      @        P       Q                   �k@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             0@        T       ]                   �c@`RI��d�?l            `e@       U       X                   �`@��FM ò?@            @Z@       V       W                   @c@`׀�:M�?,            �R@        ������������������������       �                     �?        ������������������������       �        +            @R@        Y       Z                   �s@��a�n`�?             ?@       ������������������������       �                     ;@        [       \                     P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        ,            �P@        _       �                    �?>���Rp�?�            �u@        `       y                   �b@�\����?.            �P@       a       n                   @_@#z�i��?            �D@        b       c                   `X@j���� �?             1@        ������������������������       �                     �?        d       e                    @H@      �?
             0@        ������������������������       �                     @        f       m       	          pff�?�θ�?             *@       g       h                   @]@�C��2(�?             &@        ������������������������       �                     @        i       j                    �?z�G�z�?             @        ������������������������       �                      @        k       l                    �K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        o       x                    `P@r�q��?             8@       p       u       	          033�?�C��2(�?             6@       q       r                    �?�X�<ݺ?             2@       ������������������������       �                     .@        s       t                   @p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        v       w                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        z       }                    �N@�J�4�?             9@       {       |                   �Z@�}�+r��?
             3@        ������������������������       �                     �?        ������������������������       �        	             2@        ~                          c@      �?             @        ������������������������       �                      @        �       �                   �c@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    Z@"��d`�?�            �q@        �       �                    �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �       	          pff�?vv@#_��?�            �p@        �       �                   `b@D��T��?N            �`@       �       �                    �?�S����?8            �W@       �       �                   �c@ףp=
�?.             T@       �       �                   `S@�S(��d�?+            @S@        ������������������������       �                     �?        �       �                    �?`-�I�w�?*             S@       �       �                    @L@�X�<ݺ?(             R@        ������������������������       �                     A@        �       �                    �?�KM�]�?             C@       �       �                    �?������?             1@        ������������������������       �                      @        �       �                    ]@�r����?             .@        ������������������������       �                     �?        �       �                    Y@@4և���?
             ,@        �       �                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �        
             5@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?��S���?
             .@        ������������������������       �                      @        �       �                    �F@�n_Y�K�?	             *@        ������������������������       �                     @        �       �       
             �?z�G�z�?             $@       �       �                   �r@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �F@�\��N��?             C@        ������������������������       �                     @        �       �                    �Q@����e��?            �@@       �       �                    �?f���M�?             ?@        �       �                    c@X�Cc�?             ,@        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �e@�t����?             1@       �       �                   �m@��S�ۿ?             .@       ������������������������       �                      @        �       �                   �o@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���.�6�?V            @a@       �       �                    �? _�@�Y�?F             ]@        ������������������������       �                    �C@        �       �                    �?�g<a�?3            @S@       �       �                    @J@ 7���B�?$             K@        ������������������������       �        
             0@        �       �                   �b@�}�+r��?             C@       �       �                    �J@�?�|�?            �B@        ������������������������       �                     �?        ������������������������       �                     B@        ������������������������       �                     �?        ������������������������       �                     7@        �       �                   �p@�X����?             6@       �       �                    �?�<ݚ�?             2@       �       �       	          ���@���|���?             &@        �       �                    `P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @      �?             @       �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�b�values�h)h,K ��h.��R�(KK�KK��hb�B�  !��Q��?p��1W-�?��H	9�?*�n��?�rv��?Xc"=P9�?8��18�?28��1�?�������?333333�?�������?�������?�$I�$I�?۶m۶m�?      �?                      �?�������?�������?              �?      �?      �?      �?                      �?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?              �?2�-yW��?9I�J�?s)�r)��?�����?�e˖-[�?�4iҤI�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?�����? �����?y�5���?�5��P�?�������?�������?      �?                      �?      �?        ���,d!�?8��Moz�?]t�E]�?F]t�E�?      �?      �?              �?      �?                      �?�A�A�?_�_�?      �?        I�$I�$�?۶m۶m�?              �?;�;��?;�;��?/�袋.�?F]t�E�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?5>2�ީ�?-7��X�?���)k��?��)kʚ�?9��8���?�q�q�?      �?        �������?�������?      �?                      �?{�G�z�?�z�G��?      �?              �?      �?      �?      �?      �?        UUUUUU�?�������?              �?      �?                      �?��_@�?@���?��~���?8�8��?��L��?к����?              �?      �?        �s�9��?�c�1Ƹ?      �?              �?      �?              �?      �?              �?        GX�i���?�i��F�?���>��?>����?ە�]���?�+Q��?�������?ZZZZZZ�?              �?      �?      �?              �?ى�؉��?�؉�؉�?]t�E�?F]t�E�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?�������?F]t�E�?]t�E�?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?        �z�G��?{�G�z�?�5��P�?(�����?              �?      �?              �?      �?      �?              �?      �?      �?      �?      �?                      �?              �?Y���=�?*͋?�p�?]t�E]�?F]t�E�?              �?      �?        \q�wo��?��"d
�?&���g��?���f�?^Cy�5�?(������?�������?�������?��O���?������?      �?        y�5�װ?Q^Cy��?�q�q�?��8��8�?              �?(�����?�k(���?�?xxxxxx�?      �?        �?�������?      �?        �$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�?      �?        ى�؉��?;�;��?      �?        �������?�������?�q�q�?�q�q�?              �?      �?              �?        �5��P�?y�5���?      �?        6�d�M6�?e�M6�d�?��Zk���?��RJ)��?%I�$I��?�m۶m��?              �?      �?        �?<<<<<<�?�?�������?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?              �?      �?              �?        Y�B��?���7���?�{a���?#,�4�r�?              �?�cj`?���8+�?h/�����?	�%����?              �?(�����?�5��P�?к����?*�Y7�"�?      �?                      �?      �?                      �?]t�E]�?�E]t��?�q�q�?9��8���?F]t�E�?]t�E]�?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?      �?      �?      �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�=�KhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK녔h��B�:         �                    �?�[��N�?�           ��@              Q       
             �?bz���A�?           �z@               
                    �F@4��P8O�?r            �e@                                   �?�LQ�1	�?             7@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @               	                    @��S�ۿ?             .@       ������������������������       �        
             ,@        ������������������������       �                     �?                                    �?��a_j�?b             c@                     	            �?�����	�?4            @U@        ������������������������       �                     @@                                   �?�T`�[k�?             �J@                                 `]@V������?            �B@        ������������������������       �                     "@                                  �^@��>4և�?             <@        ������������������������       �                      @                      	          ����?$��m��?             :@                                 �_@���Q��?             .@                      	          ����?�q�q�?             "@        ������������������������       �                     �?                      	             �?      �?              @        ������������������������       �                     @                                  q@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@                                  �w@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        !       .                    �?�d�K���?.            �P@        "       -       	          ����?`�Q��?             9@       #       *                    @��S���?	             .@       $       )       	          ����?�q�q�?             "@       %       &                    @K@���Q��?             @        ������������������������       �                      @        '       (                   `d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        +       ,                    �M@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        /       2                    @H@���N8�?             E@        0       1                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        3       H                    �?x�����?            �C@       4       ?                    �?�>4և��?             <@        5       6                   @`@      �?	             (@        ������������������������       �                     �?        7       8                    �K@"pc�
�?             &@        ������������������������       �                     �?        9       :                   c@ףp=
�?             $@        ������������������������       �                     @        ;       >                   �o@r�q��?             @        <       =                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        @       A                    �?      �?	             0@        ������������������������       �                     �?        B       G                   �W@��S�ۿ?             .@        C       F       	             �?      �?             @       D       E                    \@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        I       N                   �b@���!pc�?
             &@       J       M                    @      �?              @       K       L                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        O       P                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        R       u                    �?���H��?�            �o@        S       Z                    P@���}D�?*            �P@        T       U                    Z@�q�q�?             "@        ������������������������       �                      @        V       W                    �G@؇���X�?             @        ������������������������       �                     @        X       Y                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        [       d                   @\@д>��C�?#             M@        \       ]                    �E@�q�q�?
             5@        ������������������������       �                     @        ^       _                   �j@      �?             ,@        ������������������������       �                      @        `       c                   �[@�q�q�?             (@       a       b                    Z@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        e       t                    �?�L���?            �B@       f       m                    �?�#-���?            �A@        g       l                   �s@�q�q�?             @       h       k                    �I@z�G�z�?             @        i       j                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        n       o       	             �?XB���?             =@       ������������������������       �                     8@        p       q                   �d@z�G�z�?             @        ������������������������       �                     @        r       s                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        v       �                    �?�?�C+��?{             g@       w       x                    �?����?l            �d@        ������������������������       �        )             L@        y       �                   �t@d/
k�?C             [@       z       {                    @H@��-#���?B            �Z@       ������������������������       �        #            �J@        |       �                    �?�iʫ{�?            �J@        }       �                    �?����X�?             @        ~                          0c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �]@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �^@���}<S�?             G@        ������������������������       �                     1@        �       �       	            �?\-��p�?             =@       ������������������������       �                     7@        �       �                   �p@�q�q�?             @       �       �                     O@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @c@؇���X�?             5@       �       �       	          ����?      �?             (@       �       �                    �?ףp=
�?             $@        �       �                   @r@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    Z@���"�?�            0s@        �       �       	          ����?X�<ݚ�?             "@       �       �                   @X@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pe@X�����?�            �r@        �       �                   �e@����D��?8            @W@       �       �                    �M@@��,B�?6            �V@       ������������������������       �        !            �K@        �       �       	             �?������?             B@        �       �                   �[@�8��8��?             (@       ������������������������       �                     @        �       �                   �a@z�G�z�?             @        ������������������������       �                     @        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �F@�p ��?            �i@        �       �       	          hff�?�q�q�?             8@        �       �                   0p@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    b@�����H�?             2@       ������������������������       �                     0@        ������������������������       �                      @        �       �                    @R@`����e�?p            �f@       �       �                    �?��㨇,�?k            �e@       �       �                    c@`�H�/��?[             c@       �       �       
             �?Hm_!'1�?V            `b@       �       �                    @J@ =[y��?N             a@        ������������������������       �                     @@        �       �                   @i@0G���ջ?<             Z@        �       �                    ^@�θ�?             *@        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �J@x��B�R�?6            �V@        �       �                    ]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�d���?2            �U@        �       �                    �M@ףp=
�?             $@       ������������������������       �                      @        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �[@�e���@�?,            @S@        �       �                   `[@���N8�?             5@       ������������������������       �        	             *@        �       �                    �L@      �?              @        �       �       	             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     L@        �       �       	          ����?�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?      �?             @        ������������������������       �                      @        �       �       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �o@      �?             4@       �       �                    �?�q�q�?	             (@       �       �                   `@      �?              @        ������������������������       �                      @        �       �                   �b@r�q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?              @       �       �                   �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  B~�9�J�?�@c�Z�?Rh�/��?]/�ߡ�?-o�`���?iȹ�. �?Nozӛ��?d!Y�B�?      �?      �?      �?                      �?�������?�?      �?                      �?����k�?������?�?{{{{{{�?              �?"5�x+��?���!5��?o0E>��?�g�`�|�?              �?I�$I�$�?۶m۶m�?      �?        vb'vb'�?�N��N��?333333�?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?�������?333333�?              �?      �?              �?                      �?      �?      �?              �?      �?        ����?�rv��?��(\���?{�G�z�?�������?�?UUUUUU�?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��y��y�?�a�a�?UUUUUU�?UUUUUU�?      �?                      �?�A�A�?��o��o�?�m۶m��?�$I�$I�?      �?      �?      �?        F]t�E�?/�袋.�?      �?        �������?�������?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?      �?      �?        �?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?t�E]t�?F]t�E�?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �0�0�?��y��y�?&���[�?g��1��?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?a���{�?|a���?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �������?�������?�������?UUUUUU�?              �?      �?                      �?}���g�?L�Ϻ��?�A�A�?_�_�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?                      �?GX�i���?�{a���?      �?        �������?�������?      �?              �?      �?              �?      �?              �?        A�����?�5!({_�?ە�]���?,Q��+�?      �?        �Kh/���?/�����?��sH�?�琚`��?      �?        
�[���?�琚`��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        ӛ���7�?d!Y�B�?      �?        a����?�{a���?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?۶m۶m�?�$I�$I�?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �(��yھ?�Z!Ȱ$�?r�q��?�q�q�?�������?�������?      �?                      �?      �?        �3�=l}�?��DxR��?X`��?P?���O�?h�h��?`��_���?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?��+Q��?Q��+Q�?�������?�������?�������?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?      �?        X�s��C�?jc��?�'�j��?ۜ��L�?�?�������?9/���?Y�Cc�?�������?�������?              �?�؉�؉�?vb'vb'�?�؉�؉�?ى�؉��?      �?                      �?��?�����?      �?      �?      �?                      �?Ȥx�L��?�:���C�?�������?�������?              �?      �?      �?      �?                      �?�cj`?qV~B���?�a�a�?��y��y�?              �?      �?      �?�������?�������?      �?                      �?              �?              �?t�E]t�?]t�E�?      �?                      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?�������?�������?      �?      �?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?              �?      �?      �?      �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ\bshG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@0         t                    �?���-�g�?�           ��@                                 �c@�������?
           �z@                                  �Z@:�&���?.            �S@        ������������������������       �                     0@                      	          033�?��a�n`�?&             O@                                  �?^����?            �E@                                  @I@д>��C�?             =@        ������������������������       �                     &@        	       
                    [@�E��ӭ�?             2@        ������������������������       �                     @                                    P@@4և���?             ,@       ������������������������       �                     &@                                  �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                   @      �?             ,@                                  �?���|���?             &@                     	          �����X�<ݚ�?             "@        ������������������������       �                     @                                  �Z@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  �^@�KM�]�?             3@                                    O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             0@               W       
             �?V�:וd�?�            �u@               R                   pe@�^����?K            �]@               ?                   `a@�q�q�?C            @Z@       !       *                   �_@��ӭ�a�?*             R@        "       #                     F@�q�q�?             8@        ������������������������       �                      @        $       )                    @��2(&�?             6@       %       (                    �?P���Q�?             4@        &       '                   `o@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                      @        +       ,                   �`@r�q��?             H@        ������������������������       �                     @        -       >                   �`@D^��#��?            �D@       .       =                    �?D�n�3�?             C@       /       0                    �B@��S���?             >@        ������������������������       �                     @        1       8                   @d@|��?���?             ;@       2       7                   0p@p�ݯ��?             3@       3       6       	          `ff�?��S���?             .@       4       5                    �?���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        9       <       	             �?      �?              @       :       ;       
             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        @       C       
             �?<���D�?            �@@        A       B                    e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        D       O                    @��a�n`�?             ?@       E       L                   �x@ 	��p�?             =@       F       G                    �? 7���B�?             ;@       ������������������������       �                     .@        H       I       	          ����?�8��8��?             (@       ������������������������       �                     @        J       K       	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        M       N                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       Q       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       V       	          ����?@4և���?             ,@        T       U                   �e@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        X       e                    �?��F�M�?�            �l@        Y       d                   �u@��R[s�?            �A@       Z       c                    �?��X��?             <@       [       `                   0e@��H�}�?             9@       \       _                   d@��S���?             .@       ]       ^                    @H@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        a       b       	          ����?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        f       g                    �?�t�K��?{            `h@        ������������������������       �        /            �Q@        h       q                   �t@ ��+,��?L            @_@       i       j                    �I@p�,�V��?J            @^@       ������������������������       �        *            �P@        k       l                   �c@ 7���B�?              K@       ������������������������       �                    �B@        m       p                   �_@�t����?             1@        n       o                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        r       s                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        u       �                    �?������?�            0s@        v       �                    �?^H���+�?            �B@       w       �                    �?d}h���?             <@       x       }                   �b@�����?             3@       y       z                    �?؇���X�?             ,@       ������������������������       �                     $@        {       |                   `c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ~              	          `ff�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �\@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?h�WH��?�            �p@       �       �                    @ \sF��?�            @l@       �       �                    \@`2U0*��?�             l@        �       �                   �Y@      �?             8@        ������������������������       �                     �?        �       �                    @G@���}<S�?             7@        �       �                   �`@      �?              @        ������������������������       �                     @        �       �                    �F@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        �       �                   Ps@0�,���?~             i@       �       �       	          ����? }�Я��?r            @f@       �       �       	          033�?`�E���??            @X@       ������������������������       �        .            �R@        �       �                    �?�C��2(�?             6@       �       �                   �_@؇���X�?             ,@       ������������������������       �                      @        �       �                    b@�q�q�?             @       �       �                   @`@z�G�z�?             @       �       �                   �b@      �?             @        ������������������������       �                      @        �       �                    o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        3            @T@        �       �                   ``@�㙢�c�?             7@        �       �                    a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �Q@�KM�]�?
             3@       ������������������������       �        	             1@        ������������������������       �                      @        ������������������������       �                     �?        �       �                    h@�X���?             F@        �       �       	             �?�����?             5@        ������������������������       �                     &@        �       �                    �?z�G�z�?             $@        �       �                   �^@�q�q�?             @        ������������������������       �                     �?        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `@\X��t�?             7@        �       �                   `_@����X�?             @       �       �                    �?�q�q�?             @       �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          033�?     ��?             0@       ������������������������       �                     &@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  lk�w��?J��	.�?���F���?���r�.�?�o��o��?�A�A�?              �?�s�9��?�c�1��?w�qG��?�qG��?|a���?a���{�?              �?r�q��?�q�q�?      �?        �$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?]t�E]�?F]t�E�?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?(�����?�k(���?UUUUUU�?UUUUUU�?              �?      �?                      �?79ZIL�?�#����?�����?���?UUUUUU�?UUUUUU�?�8��8��?��8��8�?�������?UUUUUU�?      �?        t�E]t�?��.���?�������?ffffff�?�������?�������?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        �]�ڕ��?,Q��+�?(������?l(�����?�?�������?      �?        	�%����?{	�%���?^Cy�5�?Cy�5��?�?�������?F]t�E�?t�E]t�?              �?      �?                      �?      �?              �?      �?�������?�������?      �?                      �?              �?              �?      �?        |���?|���?      �?      �?              �?      �?        �c�1Ƹ?�s�9��?�{a���?������?h/�����?	�%����?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?      �?              �?      �?              �?      �?              �?      �?        n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?        �~]R�0�?�(�j�?X|�W|��?PuPu�?n۶m۶�?%I�$I��?{�G�z�?
ףp=
�?�������?�?ffffff�?333333�?              �?      �?                      �?�������?�������?      �?                      �?      �?              �?        �W�W�?PP�?      �?        `��"���?����Mb�?ˠT�x�?���k��?      �?        	�%����?h/�����?      �?        <<<<<<�?�?      �?      �?              �?      �?              �?              �?      �?      �?                      �?<hq��?���
�?�g�`�|�?L�Ϻ��?۶m۶m�?I�$I�$�?^Cy�5�?Q^Cy��?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?�������?�������?      �?                      �?              �?9��8���?�q�q�?              �?      �?        B{	�%��?��^B{	�?Vzja���?[X驅��?{�G�z�?���Q��?      �?      �?      �?        d!Y�B�?ӛ���7�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?g��1��?Ez�rv�?p�\��?�я~���?����??��W�?              �?F]t�E�?]t�E�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?      �?      �?                      �?              �?      �?                      �?              �?d!Y�B�?�7��Mo�?      �?      �?      �?                      �?(�����?�k(���?              �?      �?              �?        �E]t��?]t�E�?�a�a�?=��<���?              �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?!Y�B�?��Moz��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�.         l                    �?��Wޫ��?�           ��@              9                    �?$r�@&��?�            �x@                                  @E@8�����?^            �b@                                   �?      �?             D@                                   �?�eP*L��?             &@                     
             �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        	       
       	          @33�?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     =@               (       
             �?�As`�?E            �[@                      	          ����?�b��[��?"            �K@                                 �v@��
P��?            �A@                                  �?�f7�z�?             =@                     	          ����?      �?             8@        ������������������������       �                     @                                  hq@�q�q�?
             2@                                 �_@�θ�?             *@                                   �?      �?             @                                  �N@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                  �e@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                !                   �^@P���Q�?             4@        ������������������������       �                     $@        "       '                    �?ףp=
�?             $@        #       $                    �?�q�q�?             @        ������������������������       �                     �?        %       &                   ``@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        )       .                   pi@      �?#             L@        *       +                    @F@X�Cc�?	             ,@        ������������������������       �                      @        ,       -                   �h@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        /       8       	          ����?���N8�?             E@       0       7                     N@ 	��p�?             =@       1       6                    @F@h�����?             <@        2       3                   �q@�C��2(�?             &@       ������������������������       �                      @        4       5                   �r@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             1@        ������������������������       �                     �?        ������������������������       �                     *@        :       A                   �h@�Zl�i��?�            `n@        ;       @                   �^@�Fǌ��?.            �S@        <       =       
             �? �q�q�?             8@       ������������������������       �                     .@        >       ?       	             �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        #            �K@        B       C                   �Z@��
��?j            �d@        ������������������������       �                      @        D       Y       	          ����?H�ՠ&��?i            @d@        E       T       	          833�?4���C�?            �@@       F       G                    @G@ �o_��?             9@        ������������������������       �                     "@        H       I       
             �?     ��?             0@        ������������������������       �                     @        J       M                    �?�q�q�?             (@        K       L                   `^@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        N       O                    �?����X�?             @        ������������������������       �                      @        P       Q                   `m@���Q��?             @        ������������������������       �                      @        R       S                    �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        U       V                    �?      �?              @        ������������������������       �                     @        W       X       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        Z       e                    _@H*C�|F�?T             `@        [       \                   `i@      �?             8@        ������������������������       �                     �?        ]       ^                   �o@��<b���?             7@        ������������������������       �                     "@        _       d                   �\@X�Cc�?	             ,@       `       a                    �?X�<ݚ�?             "@        ������������������������       �                     @        b       c       	          ���@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        f       k                    �?@��!�Q�?D            @Z@       g       h                    �? �й���?.            @R@       ������������������������       �        #            �L@        i       j                    �Q@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        ������������������������       �                     @@        m       |                   �`@�������?�            @u@        n       w       
             �?�J���?6            @S@       o       r                    �?(L���?!            �E@        p       q                    \@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        s       v                   `X@г�wY;�?             A@        t       u                   �W@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     >@        x       y                   �V@�IєX�?             A@        ������������������������       �                     �?        z       {       	             �?Pa�	�?            �@@       ������������������������       �                     @@        ������������������������       �                     �?        }       �                    �K@J���?�            pp@       ~       �       
             �?�ˈ��@�?x            �h@               �                    @�����?            �L@       �       �                    �G@ \� ���?            �H@        �       �                   �[@P���Q�?             4@        ������������������������       �                     �?        ������������������������       �        
             3@        �       �                   �b@����"�?             =@       �       �       	          ����? �o_��?             9@       �       �                   �\@r�q��?             2@        �       �                   `d@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �b@@4և���?	             ,@        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   0a@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �r@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        Y            �a@        �       �                   �a@      �?$            �P@        ������������������������       �                     @        �       �                    �?�G�z��?!             N@       �       �                     O@z�G�z�?             >@       �       �                    �?�C��2(�?
             6@        �       �                   (s@����X�?             @       �       �                   8p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     .@        �       �                    b@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                    �P@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �q@�z�G��?             >@       �       �                    �?և���X�?             5@        �       �                   �b@X�<ݚ�?             "@       �       �                   0b@r�q��?             @        ������������������������       �                     @        �       �       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                     M@      �?             @        ������������������������       �                     �?        �       �                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �N@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B�  +^�ɑA�?�P47��?�լ?��?���0�?��{���?�B���?      �?      �?]t�E�?t�E]t�?�$I�$I�?�m۶m��?              �?      �?              �?      �?      �?                      �?              �?�9	ą��?���w���?־a��?� O	��?PuPu�?_�_��?a���{�?O#,�4��?      �?      �?              �?UUUUUU�?UUUUUU�?ى�؉��?�؉�؉�?      �?      �?      �?      �?      �?                      �?              �?      �?        �������?333333�?              �?      �?                      �?      �?        �������?ffffff�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?      �?%I�$I��?�m۶m��?              �?      �?      �?      �?                      �?��y��y�?�a�a�?������?�{a���?�m۶m��?�$I�$I�?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �����H�?�"e����?�3���?1���M��?UUUUUU�?�������?              �?�q�q�?�q�q�?              �?      �?                      �?�18���?��18��?      �?        {	�%���?������?'�l��&�?m��&�l�?�Q����?
ףp=
�?              �?      �?      �?              �?�������?�������?�������?333333�?      �?                      �?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�!oȫ?�7�yC�?      �?      �?      �?        ��Moz��?��,d!�?              �?�m۶m��?%I�$I��?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?8�8��? �����?����?����Ǐ�?              �?      �?      �?              �?      �?                      �?�������?�������?qV~B���?����15�?w�qG��?⎸#��?r�q��?�q�q�?              �?      �?        �?�?      �?      �?              �?      �?                      �?�?�?              �?|���?|���?      �?                      �?�m�o��?��K>@��?T��~�?\e
�d�?Q^Cy��?^Cy�5�?
^N��)�?և���X�?ffffff�?�������?              �?      �?        	�=����?�i��F�?
ףp=
�?�Q����?�������?UUUUUU�?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?                      �?      �?      �?              �?      �?              �?              �?      �?      �?        �������?�������?�������?�������?F]t�E�?]t�E�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?ffffff�?333333�?�$I�$I�?۶m۶m�?�q�q�?r�q��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJj�c;hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKᅔh��B@8         h                   �`@$~��,��?�           ��@               E       	          ����?�`��9�?�            �u@                                   �?,z�?���?t            �f@                                  �?�E���?@            @X@        ������������������������       �                     9@                                  �\@      �?2             R@               
       
             �?�t����?             A@              	       
             �?�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@                                   [@"pc�
�?             &@                     	          @33�?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?                                  `]@�����?             C@        ������������������������       �                      @                                   �?�E��ӭ�?             B@                                  �? �Cc}�?             <@                      
             �?և���X�?             @                                 �`@���Q��?             @                     	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             5@                                  �`@      �?              @        ������������������������       �                     @                                   b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        !       :       
             �?؇���X�?4             U@       "       %                    �?����1�?,            @R@        #       $                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        &       /                    l@t�e�í�?(            �P@       '       (                   pi@`Ql�R�?            �G@       ������������������������       �                     B@        )       .                    �?�C��2(�?             &@       *       +                    �?      �?              @       ������������������������       �                     @        ,       -                   @\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        0       1                   �l@z�G�z�?             4@        ������������������������       �                     �?        2       9                    �?�S����?             3@       3       4                    _@�IєX�?             1@        ������������������������       �                      @        5       8                   xp@�����H�?             "@        6       7                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ;       <                    Z@�eP*L��?             &@        ������������������������       �                      @        =       B                    �?X�<ݚ�?             "@       >       ?       	          ����?�q�q�?             @        ������������������������       �                     @        @       A                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        C       D                   @b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        F       O                   `\@��O���?k            @e@        G       H                    �?�n_Y�K�?             *@        ������������������������       �                      @        I       J                    �?���!pc�?             &@        ������������������������       �                     �?        K       L       
             �?z�G�z�?             $@        ������������������������       �                     @        M       N                    �K@      �?             @       ������������������������       �                      @        ������������������������       �                      @        P       Y                    �?�E����?d            �c@        Q       R                    @O@      �?             <@       ������������������������       �                     1@        S       T                   �`@���|���?             &@        ������������������������       �                     @        U       V                   pb@      �?              @        ������������������������       �                     @        W       X                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        Z       _                     E@0Ƭ!sĮ?Q             `@        [       ^                    `@���Q��?             @        \       ]       	             @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        `       c                   @^@0�z��?�?M             _@        a       b                   ``@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        d       e                   P`@@���a��?E            �\@       ������������������������       �        ?            @Z@        f       g                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        i       �                    �?6R��P��?�            �w@        j       �       	          ����?b����?V            �_@       k       x                   �i@(ǯt��?3            �R@        l       w                    �?��2(&�?             6@       m       n       
             �?     ��?             0@        ������������������������       �                      @        o       v                    �L@      �?              @       p       q                    �?���Q��?             @        ������������������������       �                     �?        r       u                   @`@      �?             @        s       t                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        y       z                   �a@�	j*D�?"             J@        ������������������������       �                     ,@        {       �       
             �?D�n�3�?             C@        |                           �?X�<ݚ�?             "@       }       ~                    @L@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                     F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�f7�z�?             =@       �       �                   0e@�d�����?             3@       �       �                    �E@X�<ݚ�?	             "@        ������������������������       �                      @        �       �                    �?����X�?             @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �d@�z�G��?             $@       �       �                   @c@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   e@4��?�?#             J@       �       �                    �? �q�q�?              H@        �       �                   pc@8�Z$���?
             *@       ������������������������       �                     $@        �       �                     G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �A@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��-���?�            p@        �       �                    �K@��y� �?;            @W@       �       �       
             �? �й���?/            @R@        �       �                   �b@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �        "            �J@        �       �                   �e@��Q��?             4@       �       �                    �?�r����?             .@       �       �                   �b@�8��8��?	             (@        �       �                    @N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �K@���01m�?a            �d@       �       �       
             �?>A�F<�?D            �\@        �       �                    �?��J�fj�?            �B@        ������������������������       �                     @        �       �                   �r@�4�����?             ?@       �       �                     G@���B���?             :@        �       �       	          ����?���|���?             &@        ������������������������       �                     @        �       �                   �o@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    b@��S�ۿ?             .@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �        /            @S@        �       �                   m@���Q��?             I@       �       �                   �^@�q�q�?             8@        ������������������������       �                      @        �       �                    �?���|���?             6@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             2@       �       �                   �b@և���X�?	             ,@        ������������������������       �                     @        �       �                    �?���!pc�?             &@       �       �                   0l@؇���X�?             @       ������������������������       �                     @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?�θ�?             :@       �       �                    b@�X�<ݺ?             2@       ������������������������       �                     .@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   Ps@      �?              @       �       �                    �?r�q��?             @       �       �                   p`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  ��C�l��??+^�ɑ�?���X:�?-~�����?�.�^���?�h�P�?tT����?W?���?      �?              �?      �?�������?�������?d!Y�B�?�Mozӛ�?      �?                      �?/�袋.�?F]t�E�?�������?�������?      �?                      �?              �?Q^Cy��?^Cy�5�?              �?�q�q�?r�q��?%I�$I��?۶m۶m�?�$I�$I�?۶m۶m�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?Ĉ#F��?�Ν;w��?UUUUUU�?UUUUUU�?      �?                      �?�rv��?�1����?W�+�ɕ?}g���Q�?              �?F]t�E�?]t�E�?      �?      �?              �?      �?      �?      �?                      �?              �?�������?�������?      �?        ^Cy�5�?(������?�?�?              �?�q�q�?�q�q�?      �?      �?      �?                      �?              �?      �?        ]t�E�?t�E]t�?              �?r�q��?�q�q�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?�������?ى�؉��?;�;��?      �?        t�E]t�?F]t�E�?      �?        �������?�������?              �?      �?      �?              �?      �?        �����?�}��	��?      �?      �?              �?]t�E]�?F]t�E�?      �?              �?      �?              �?�������?�������?      �?                      �?����?����?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�B!��?|���{�?�q�q�?�q�q�?              �?      �?        ���ρ?�uI�ø�?              �?�������?�������?              �?      �?        Z�In%8�?M�l#���?�eY�eY�?5M�4M��?���g��?S�n0E�?t�E]t�?��.���?      �?      �?              �?      �?      �?333333�?�������?              �?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?vb'vb'�?;�;��?      �?        l(�����?(������?r�q��?�q�q�?�$I�$I�?۶m۶m�?              �?      �?              �?      �?              �?      �?        O#,�4��?a���{�?Cy�5��?y�5���?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?        333333�?ffffff�?      �?      �?              �?      �?              �?        ى�؉��?�N��N��?UUUUUU�?�������?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?Y�X�X��?�b�b�b�??���O?�?X`��?����Ǐ�?����?ffffff�?�������?      �?                      �?      �?        �������?ffffff�?�������?�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?                      �?���|�?�cp>��?������?Cy�5��?к����?�"�u�)�?      �?        ��RJ)��?���Zk��?ى�؉��?��؉���?F]t�E�?]t�E]�?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�������?      �?      �?              �?      �?                      �?      �?              �?        �������?333333�?�������?�������?              �?]t�E]�?F]t�E�?      �?        r�q��?�q�q�?۶m۶m�?�$I�$I�?      �?        t�E]t�?F]t�E�?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?      �?      �?                      �?      �?        �؉�؉�?ى�؉��?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJGԙGhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKŅ�h��B@1         |       
             �?�/�$�y�?�           ��@              !                    �?$�P�Gn�?            {@                                   �?��
ц��?+            @P@                                  b@">�֕�?            �A@                                 �\@      �?             6@        ������������������������       �                     @                                  �r@b�2�tk�?             2@                                  a@����X�?
             ,@       	       
       	          pff�?r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @                                  hu@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@                      	          ����?z�G�z�?             >@                                   Z@����X�?             @        ������������������������       �                      @                                  �k@���Q��?             @        ������������������������       �                     �?                                  p@      �?             @        ������������������������       �                      @                                  �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                       	          `ff�?�nkK�?             7@                      	          ����?؇���X�?             @        ������������������������       �                     @                                  �_@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     0@        "       S                   �a@�d�W��?�            w@       #       L                    `P@���۟�?�            `q@       $       )       
             �?��a��?�            @n@        %       (                    �?�+$�jP�?             ;@        &       '                   @`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        *       5                   �[@�V���?�            �j@        +       4                    �L@�S����?             3@        ,       3                    �?���!pc�?             &@       -       .                   @Z@      �?              @        ������������������������       �                     �?        /       2                    �K@և���X�?             @       0       1                   �m@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        6       E       	          ����?`�(c�?v            �h@        7       8       	          ����?0��P�?3            �T@       ������������������������       �                    �G@        9       :                   Pn@؇���X�?            �A@       ������������������������       �                     6@        ;       D                   `@�n_Y�K�?	             *@       <       =                    Z@���!pc�?             &@        ������������������������       �                     @        >       C                    �?և���X�?             @       ?       @                    @N@z�G�z�?             @        ������������������������       �                     @        A       B                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        F       K                    �J@�Ru߬Α?C            �\@        G       J                   �_@�Ń��̧?             E@        H       I                   �^@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �        +             R@        M       R                    �?r�q��?             B@        N       Q                   @p@�q�q�?             "@       O       P       	          ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ;@        T       U                   �Z@����X�?9            �V@        ������������������������       �                     @        V       c                    �?�/,Tg�?7             U@        W       X                    @L@��p\�?            �D@       ������������������������       �                     6@        Y       b                   �a@�S����?             3@       Z       a                   �q@���!pc�?             &@       [       \                   @`@      �?             @        ������������������������       �                     �?        ]       `                     P@���Q��?             @       ^       _                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        d       u                   �n@�lg����?            �E@       e       p                   �`@      �?             :@       f       o       	          `ff@�t����?             1@       g       h                   �\@؇���X�?	             ,@        ������������������������       �                     �?        i       j                    @L@$�q-�?             *@       ������������������������       �                      @        k       n       	          ����?z�G�z�?             @       l       m                    �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        q       r                   pk@�����H�?             "@       ������������������������       �                     @        s       t                    @O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        v       {                   f@@�0�!��?             1@       w       z                    @K@��S�ۿ?
             .@        x       y                   0c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        }       �                    �?��J��?�            �r@        ~                          d@=QcG��?;            �W@       ������������������������       �        "            �I@        �       �                   @d@(L���?            �E@        ������������������������       �                     @        �       �                   �Z@��(\���?             D@        �       �                   �X@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?г�wY;�?             A@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @@        �       �       	            �?�C;���?�            �i@       �       �                    @M@L�
�$�?_            �a@       �       �                    �?�S���?R             ^@       �       �                   @E@h�����?N             \@        �       �                    �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @L@�O4R���?I            �Z@       ������������������������       �        B            @X@        �       �                   �l@�<ݚ�?             "@       ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �I@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �P@�G��l��?             5@       �       �                    �?X�<ݚ�?
             2@        �       �                    �?����X�?             @       �       �                   @_@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    b@���!pc�?             &@       �       �       	          ����?���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    ]@�G\�c�?&            @P@        ������������������������       �                     @        �       �                   `_@��o	��?$             M@        ������������������������       �                     "@        �       �                    �?Tt�ó��?            �H@       �       �       	             @�q�q�?             B@       �       �                    �J@��a�n`�?             ?@        �       �                   0`@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @`@���}<S�?             7@        �       �                   `k@�<ݚ�?             "@        ������������������������       �                     @        �       �       	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             ,@        ������������������������       �                     @        �       �                   p`@�θ�?             *@        ������������������������       �                      @        �       �                   `W@�C��2(�?	             &@        �       �       	             �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  L�f���?Z�L��?��_ǯ��?P(�?�;�;�?�؉�؉�?�A�A�?_�_��?      �?      �?              �?�8��8��?9��8���?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?                      �?�������?�������?�$I�$I�?�m۶m��?              �?�������?333333�?      �?              �?      �?              �?      �?      �?              �?      �?        �Mozӛ�?d!Y�B�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?        ?uG���?X�j��?����j�?��a����?���|���?��2(&�?B{	�%��?/�����?�������?UUUUUU�?      �?                      �?              �?��V!�n�?D��=��?^Cy�5�?(������?t�E]t�?F]t�E�?      �?      �?              �?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?                      �?              �?և���X�?��)x9�?8��18�?���|�?              �?�$I�$I�?۶m۶m�?              �?ى�؉��?;�;��?t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?      �?      �?                      �?      �?              �?        p�}��?���#��?�a�a�?��<��<�?�?�������?              �?      �?                      �?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?              �?�$I�$I�?�m۶m��?      �?        =��<���?1�0��?��+Q��?�]�ڕ��?              �?^Cy�5�?(������?t�E]t�?F]t�E�?      �?      �?              �?333333�?�������?      �?      �?      �?                      �?              �?              �?              �?�}A_��?}A_��?      �?      �?�������?�������?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�q�q�?�q�q�?              �?      �?      �?              �?      �?        �������?ZZZZZZ�?�?�������?�������?�������?      �?                      �?              �?      �?        ~��K~�?:m���?x6�;��?AL� &W�?      �?        ⎸#��?w�qG��?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?        �?�?      �?      �?              �?      �?              �?        a����t�?>�Tr^�?qJ��O$�?{�e�ݾ?""""""�?�����ݭ?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?        :�&oe�?�x+�R�?      �?        9��8���?�q�q�?      �?              �?      �?              �?      �?              �?      �?      �?                      �?1�0��?��y��y�?�q�q�?r�q��?�m۶m��?�$I�$I�?333333�?�������?              �?      �?              �?        t�E]t�?F]t�E�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        [��Z���?S+�R+��?              �?������?���{�?              �?h�����?/�����?UUUUUU�?UUUUUU�?�c�1��?�s�9��?      �?      �?              �?      �?        ӛ���7�?d!Y�B�?9��8���?�q�q�?      �?              �?      �?              �?      �?              �?                      �?�؉�؉�?ى�؉��?      �?        F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��AhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@/         p                    �?z��K���?�           ��@              3                    �?1`�N�?�            y@               *                    �?z�):���?X            �b@              )       	          ���@�s��:��?D            �\@                     
             �?�	#i���??            �Z@                      	          ����?p�v>��?            �G@        ������������������������       �                     4@                                  �a@|��?���?             ;@       	                           �?���|���?             6@        
              	          ����?����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                  �^@z�G�z�?             .@                                  �F@      �?              @        ������������������������       �                     @                                  �^@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   T@���*�?#             N@                      	          @33�?���Q��?             @        ������������������������       �                     �?                                   a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �b@t�6Z���?            �K@       ������������������������       �                     :@               $                    �L@�c�Α�?             =@              #                    ^@�㙢�c�?             7@               "                    q@���|���?             &@               !                     E@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        %       &                   �o@�q�q�?             @        ������������������������       �                      @        '       (                   �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        +       0                    l@r�q��?             B@       ,       /                    �?(;L]n�?             >@        -       .                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     <@        1       2       
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        4       [       
             �?���+[��?�            `o@       5       P       	          ����?�
���x�?�             k@        6       C                    �?� y���?,            �P@       7       <                    �? i���t�?             �H@        8       9                    �?������?             .@        ������������������������       �                     @        :       ;                   �s@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        =       >       
             �?г�wY;�?             A@        ������������������������       �                      @        ?       B                   �[@      �?             @@        @       A                   @[@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     3@        D       E                    �?�q�q�?             2@        ������������������������       �                      @        F       G       	             �?      �?
             0@        ������������������������       �                     @        H       O                     M@���Q��?             $@       I       J                   @\@      �?              @        ������������������������       �                     @        K       N                    b@z�G�z�?             @       L       M                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Q       R                   �b@��
���?\            �b@       ������������������������       �        A             Z@        S       T                     F@���}<S�?             G@        ������������������������       �                      @        U       Z                   �\@���7�?             F@        V       Y       	             @�KM�]�?             3@       W       X                   �[@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     9@        \       i                   �a@ҳ�wY;�?             A@       ]       ^                    �?�q�q�?             8@        ������������������������       �                     �?        _       d       	          ����?�㙢�c�?             7@        `       c                   �d@�q�q�?             "@       a       b                   �a@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        e       h                   `U@@4և���?
             ,@       f       g       	          `ff�?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        j       m                    n@�z�G��?             $@       k       l                    �N@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        n       o                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        q       �       
             �?Ɨ�v2U�?�            �t@        r       �       	          ����?�R�G�?K            @_@        s       �                   �b@tk~X��?             B@       t       w                    �?������?             ;@        u       v                    e@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        x                          �[@�X�<ݺ?             2@        y       ~                    �?�����H�?             "@       z       }                    �?      �?             @        {       |                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     "@        �       �                    �?���R��?5            @V@        �       �       	          ����?�����?             3@        ������������������������       �                      @        �       �                    �?������?             1@        ������������������������       �                     @        �       �                   �\@�q�q�?
             (@        ������������������������       �                     @        �       �                   Xq@      �?              @       �       �                   �j@�q�q�?             @        ������������������������       �                     �?        �       �                    �K@z�G�z�?             @        ������������������������       �                      @        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?���Q��?%            �Q@        �       �                    o@�r����?             .@       ������������������������       �                     &@        �       �                    �M@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   P`@���!pc�?            �K@       �       �       	             �?\�Uo��?             C@        ������������������������       �                     @        �       �                   �a@     ��?             @@        ������������������������       �                     $@        �       �       	          `ff@8�A�0��?	             6@       �       �       	          `ff�?�q�q�?             (@       �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �\@z�G�z�?             $@        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@        �       �                    �O@ ��WV�?�             j@       �       �                   Pc@��Μ�V�?y             h@        �       �       	            �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     L@��K2��?u            �g@       ������������������������       �        h             e@        �       �                   0b@�KM�]�?             3@        �       �       	          @33�?����X�?             @       ������������������������       �                     @        �       �                    q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        �       �                    �?�q�q�?             .@        ������������������������       �                      @        �       �                   p@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  K�ۚ��?�)|�� �?��N���?�{^��V�?q=
ףp�?H�z�G�?��k(��?�k(���?|d�S��?7��XQ�?L� &W�?ڨ�l�w�?              �?{	�%���?	�%����?]t�E]�?F]t�E�?�$I�$I�?�m۶m��?      �?                      �?�������?�������?      �?      �?      �?        �������?333333�?              �?      �?              �?                      �?""""""�?wwwwww�?�������?333333�?      �?              �?      �?              �?      �?        X���oX�?��)A��?      �?        5�rO#,�?�{a���?�7��Mo�?d!Y�B�?]t�E]�?F]t�E�?9��8���?�q�q�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?UUUUUU�?�������?�?�������?      �?      �?              �?      �?                      �?�������?UUUUUU�?              �?      �?        �';r���?���Ɏ�?��Fd#��?�&w����?~5&��?z�rv��?����X�?/�����?�?wwwwww�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?�?              �?      �?      �?;�;��?�؉�؉�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?�������?333333�?      �?      �?      �?        �������?�������?      �?      �?              �?      �?                      �?              �?O贁N�?&�X�%�?              �?d!Y�B�?ӛ���7�?      �?        F]t�E�?�.�袋�?(�����?�k(���?UUUUUU�?�������?              �?      �?                      �?              �?�������?�������?�������?UUUUUU�?      �?        d!Y�B�?�7��Mo�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?      �?        �$I�$I�?n۶m۶�?�$I�$I�?۶m۶m�?              �?      �?                      �?ffffff�?333333�?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        O}Q����?b]#V�?�~j�t��?��ʡE��?9��8���?r�q��?{	�%���?B{	�%��?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?��8��8�?�q�q�?�q�q�?      �?      �?      �?      �?      �?                      �?              �?              �?              �?              �?ؽ�u�{�?�E(B�?Q^Cy��?^Cy�5�?              �?xxxxxx�?�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?333333�?�������?�?      �?              �?      �?      �?                      �?t�E]t�?F]t�E�?6��P^C�?�5��P^�?      �?              �?      �?              �?/�袋.�?颋.���?�������?�������?      �?      �?              �?      �?      �?              �?      �?              �?        �������?�������?�������?333333�?              �?      �?                      �?              �?O��N���?;�;��?�GJȩ��?�n�Տ?�������?�������?      �?                      �?��Q�٨�?W�+�Ʌ?      �?        �k(���?(�����?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?�m۶m��?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ,�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKͅ�h��B@3         x       
             �?8}�ý�?�           ��@              a                    �?:_q�q�?
           �z@                                   �?���h���?�            s@                                   �D@���h%��?'            �O@        ������������������������       �                     @                                  @[@6�iL�?$            �M@        ������������������������       �                     @                                  d@4և����?"             L@       	              	             @���j��?             G@       
                          �c@8�Z$���?            �C@                                  �?d}h���?             <@                                  �N@�t����?             1@                                 Pc@"pc�
�?             &@                                  �K@ףp=
�?             $@       ������������������������       �                     @                                  @`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                    K@���|���?	             &@        ������������������������       �                     @                                   d@�q�q�?             @                     	          033�?z�G�z�?             @                                  `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     $@        !       ^       	          `ff@��2(&�?�            @n@       "       C                    �?H�f�i��?�            @m@       #       2                    �?�8��?f            �d@        $       )                   �k@�������?             A@        %       (                    `@@4և���?
             ,@        &       '                   �^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        *       +       	          ����?���Q��?             4@        ������������������������       �                     "@        ,       /                    @H@���!pc�?             &@        -       .                    �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        0       1       	          033�?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        3       4                   �Z@pJQg���?O            �`@        ������������������������       �                     �?        5       <       	          033@����e��?N            �`@       6       ;                   �i@@���a��?@            �\@        7       8                    �?г�wY;�?             A@       ������������������������       �                     >@        9       :       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        +            @T@        =       B                    `@�IєX�?             1@        >       A       	          ���@z�G�z�?             @        ?       @                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             (@        D       E       
             �?.��<�?(            �P@        ������������������������       �                     @        F       I                     E@     ��?%             P@        G       H                    �A@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        J       Y                    �O@�S����?            �L@       K       T                    �?ףp=
�?             I@       L       S                     N@      �?             @@       M       R                   �`@z�G�z�?             4@       N       O                     I@���Q��?             $@        ������������������������       �                     @        P       Q                   �b@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     (@        U       V                   �`@�X�<ݺ?	             2@       ������������������������       �                     "@        W       X                    �M@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        Z       [       	          ����?և���X�?             @        ������������������������       �                     @        \       ]                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        _       `                   �c@      �?              @       ������������������������       �                     @        ������������������������       �                     @        b       u                   �r@\����?Q            @^@       c       d                    �?���7�?J            �[@       ������������������������       �        8            �U@        e       n                    �?��<b���?             7@        f       g                   �\@      �?              @        ������������������������       �                     �?        h       m                   �n@����X�?             @       i       j                   @_@      �?             @        ������������������������       �                     �?        k       l                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        o       t       	          `ff@�r����?
             .@       p       q                    �?@4և���?	             ,@       ������������������������       �                     $@        r       s                   �_@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        v       w                   t@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        y       �                   �S@�������?�            @s@        z       �                   �_@:ɨ��?            �@@        {       �       	          ����?@�0�!��?	             1@        |                           �?և���X�?             @       }       ~                   �c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?     ��?             0@       �       �                   `]@�q�q�?             "@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�@�' �?�            0q@       �       �                   pc@�A6��Ľ?�            @n@       �       �                   �p@ g�yB�?Q             `@       ������������������������       �        ?            �Z@        �       �                   �p@���}<S�?             7@        ������������������������       �                     �?        �       �       	          ����?���7�?             6@       �       �                    �?�IєX�?             1@        �       �                    @L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     @        �       �                    �?��(�?H            @\@        �       �                    �?�û��|�?             7@        �       �       	             �?���!pc�?             &@       �       �                   �r@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?	             (@        ������������������������       �                     �?        �       �       	          ����?�eP*L��?             &@       �       �                    �G@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �d@`Ӹ����?9            �V@        �       �                    �?<���D�?            �@@        ������������������������       �                      @        �       �                   xt@�J�4�?             9@       �       �                    c@      �?             8@       �       �                    d@�X�<ݺ?             2@       ������������������������       �                     (@        �       �                     @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        (            �L@        �       �                    �?���|���?            �@@       �       �       	          ����?�c�Α�?             =@        �       �                    �Q@և���X�?
             ,@       �       �                    �?�q�q�?	             (@        ������������������������       �                     �?        �       �                   @`@���|���?             &@        �       �                   �q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?؇���X�?             @        ������������������������       �                      @        �       �                    h@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B�  a[ӿc�?PR Np�?��PI7��?Yޫ-r��?pk�$��?$����?v]�u]��?EQEQ�?              �?ylE�pR�?'u_[�?              �?%I�$I��?n۶m۶�?ozӛ���?!Y�B�?;�;��?;�;��?I�$I�$�?۶m۶m�?<<<<<<�?�?/�袋.�?F]t�E�?�������?�������?      �?              �?      �?              �?      �?                      �?      �?        ]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?                      �?      �?        t�E]t�?��.���?�������?�����?7Āt,e�?y�oqZ��?�������?�������?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?�������?333333�?              �?F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�qA��?s���7G�?      �?        |���?�>����?���ρ?�uI�ø�?�?�?              �?      �?      �?              �?      �?                      �?�?�?�������?�������?      �?      �?              �?      �?                      �?              �?o�Wc"=�?IT�n��?      �?              �?      �?�m۶m��?�$I�$I�?              �?      �?        ^Cy�5�?(������?�������?�������?      �?      �?�������?�������?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�q�q�?��8��8�?              �?�q�q�?�q�q�?              �?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?      �?      �?              �?      �?        "pc�
�?���|���?F]t�E�?�.�袋�?              �?��Moz��?��,d!�?      �?      �?      �?        �$I�$I�?�m۶m��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�?�������?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?              �?        F]t�E�?]t�E]�?      �?                      �?{�����?�����?e�M6�d�?N6�d�M�?�������?ZZZZZZ�?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�{�����?����?��Z=;�?�eP*L��?�����?����?      �?        ӛ���7�?d!Y�B�?              �?�.�袋�?F]t�E�?�?�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �Ź�Q�?�8�1�s�?8��Moz�?��,d!�?F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?        ]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?        ?�>��?l�l��?|���?|���?      �?        �z�G��?{�G�z�?      �?      �?��8��8�?�q�q�?      �?        �������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        F]t�E�?]t�E]�?�{a���?5�rO#,�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?        ]t�E]�?F]t�E�?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?                      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJf��'hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKŅ�h��B@1         �       
             �?�3u���?�           ��@              I                    �?����؜�?           pz@                                  `\@֭��F?�?r            �g@                                   �? 7���B�?             ;@       ������������������������       �                     4@                                  `X@؇���X�?             @               
                    �?�q�q�?             @              	                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               &                    �?�h��?[             d@                                  �k@.��<�?&            �P@                                  �?�?�|�?            �B@                                    H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     A@                                  �^@��S���?             >@                                   �?z�G�z�?             .@        ������������������������       �                     @                                   @D@      �?              @        ������������������������       �                     �?                                  �Z@����X�?             @        ������������������������       �                     �?                                  �^@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @               %                    �?������?
             .@              $                    �M@8�Z$���?	             *@                !                   �`@����X�?             @        ������������������������       �                     @        "       #                   b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        '       F                    �?�[�IJ�?5            �W@       (       1                    �?�G�z��?/             T@        )       0                    �?�חF�P�?             ?@       *       /                   `c@ܷ��?��?             =@       +       .                   �b@ 7���B�?             ;@        ,       -                   �b@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                      @        ������������������������       �                      @        2       3                    @B@�`���?            �H@        ������������������������       �                     @        4       5                    ]@�D����?             E@        ������������������������       �                     @        6       A                   �b@4�B��?            �B@       7       :       	             �?����"�?             =@       8       9                   @a@�t����?
             1@        ������������������������       �                      @        ������������������������       �                     .@        ;       @                   d@      �?             (@       <       =                    �N@"pc�
�?             &@       ������������������������       �                      @        >       ?                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        B       C                   pq@      �?              @       ������������������������       �                     @        D       E                   e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        G       H                   @`@d}h���?             ,@        ������������������������       �                     @        ������������������������       �                     &@        J       �                    �N@8���@�?�            `m@       K       Z                    �?�j��b�?~             f@        L       Y                   �b@8����?             7@       M       V                    �?���N8�?             5@       N       Q                    _@@�0�!��?             1@        O       P                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        R       S                    @L@�r����?             .@       ������������������������       �                     (@        T       U       	          `ff�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        W       X                   �o@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        [       ~                    c@@4և���?m            @c@       \       ]                   �Z@�c!�^�?i            @b@        ������������������������       �                     �?        ^       c                   @X@����=O�?h             b@        _       b                   l@      �?              @        `       a                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        d       e                    �?���Z�?b             a@        ������������������������       �                     D@        f       {                   �s@h�a��?I            @X@       g       z                   �o@`Ӹ����?B            �V@       h       w                    @N@p��%���?3            @Q@       i       v                   �l@���7�?0            �P@       j       u                   pl@�1�`jg�?(            �K@       k       l       	          033�? 7���B�?'             K@        ������������������������       �                     8@        m       p                   �`@��S�ۿ?             >@       n       o                    \@ ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        q       r                    �?      �?             @        ������������������������       �                      @        s       t                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        x       y                   `^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        |       }       	          ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @               �                     M@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    \@ _�@�Y�?&             M@        �       �                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        $            �K@        �       �                   @E@v�9ч.�?�            ps@        �       �                    �?���"͏�?            �B@        �       �                     E@      �?
             0@        ������������������������       �                      @        �       �       	            �?����X�?	             ,@        ������������������������       �                     @        �       �                     P@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                   �_@؇���X�?             5@        ������������������������       �                     "@        �       �                    �?      �?             (@       �       �                    @K@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?`cjg�?�             q@       �       �                    �?���X=P�?�            �n@        �       �                   �a@z�G�z�?'            �K@        ������������������������       �                     >@        �       �                    �M@� �	��?             9@       �       �       	          ����?�q�q�?             5@       �       �                    @F@     ��?             0@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �`@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             @��s��?w            �g@       �       �                   �c@@>ZAɥ�?u            `g@       �       �                    �?����X�?D             \@       �       �                     L@     ��?'             P@       ������������������������       �        !             M@        �       �                    p@r�q��?             @        ������������������������       �                     @        �       �                     M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     H@        �       �                    @M@Х-��ٹ?1            �R@       ������������������������       �        -             Q@        �       �                   @b@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?l��[B��?             =@       �       �                   `u@�z�G��?             4@       �       �                    �L@�<ݚ�?             2@        �       �                    �H@      �?              @        ������������������������       �                     @        �       �                   Pe@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �d@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  k�w죻�?��	."�?Q�oa��?�k���?br1���?�F}g���?h/�����?	�%����?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?�.>9�?��h�`��?o�Wc"=�?IT�n��?к����?*�Y7�"�?UUUUUU�?UUUUUU�?              �?      �?                      �?�?�������?�������?�������?      �?              �?      �?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?        �?wwwwww�?;�;��?;�;��?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?                      �?      �?        ���
b�?m�w6�;�?ffffff�?333333�?�Zk����?��RJ)��?��=���?a���{�?	�%����?h/�����?�q�q�?�q�q�?      �?                      �?      �?                      �?              �?����S�?և���X�?              �?�0�0�?z��y���?              �?�Y7�"��?L�Ϻ��?	�=����?�i��F�?<<<<<<�?�?              �?      �?              �?      �?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?              �?      �?              �?      �?        ۶m۶m�?I�$I�$�?      �?                      �? ��§��?�"��i�?��/���?�N��?8��Moz�?d!Y�B�?��y��y�?�a�a�?�������?ZZZZZZ�?      �?      �?              �?      �?        �?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?        �$I�$I�?n۶m۶�?Ĉ#F��?t�Ν;w�?      �?        ��RA�/�?U��K��?      �?      �?      �?      �?              �?      �?                      �?T{N���?�J���?              �?���Id�?�D�a�Y�?l�l��??�>��?ہ�v`��?�g��%�?F]t�E�?�.�袋�?�־a�?A��)A�?h/�����?	�%����?              �?�?�������?;�;��?O��N���?      �?                      �?      �?      �?              �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?              �?      �?        �{a���?#,�4�r�?UUUUUU�?UUUUUU�?      �?                      �?              �?<�5��?ϣ�)�?*�Y7�"�?v�)�Y7�?      �?      �?      �?        �$I�$I�?�m۶m��?      �?        F]t�E�?]t�E�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?���L_%�?�J�վ?�j򸳄�?]�l8bڳ?�������?�������?      �?        �Q����?)\���(�?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?              �?        �������?�������?              �?      �?                      �?q�����?�X�0Ҏ�?%��j�$�?a�2a�?n۶m۶�?�$I�$I�?     ��?      �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        K~��K�?O贁N�?      �?        ۶m۶m�?�$I�$I�?              �?      �?                      �?���=��?GX�i���?333333�?ffffff�?�q�q�?9��8���?      �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?�������?�������?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJy"rhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�/         �       
             �?�$���?�           ��@              =                   a@ lee�i�?           �z@              :                    �R@P�Q���?�            �p@                                  �?�U�=���?�            �p@                                  0l@R�}e�.�?             :@        ������������������������       �                     *@               
       	          ����?��
ц��?
             *@              	                    w@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                      
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @               9                    �?8Z��Up�?�            �m@              8                   `@`ۘV�?p            @e@              )                    `@������?b             b@               &       	          033@��k=.��?             �G@              %       	          `ff�?(L���?            �E@              "                    �?�+e�X�?             9@                                 �^@"pc�
�?             6@                                  �?�KM�]�?             3@        ������������������������       �                     @                                  `Z@r�q��?             (@                                  X@����X�?             @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                     �?                                   @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                !                    Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        #       $                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             2@        '       (                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        *       +                    �D@@9G��?B            �X@        ������������������������       �                      @        ,       -                   `[@@��8��?A             X@        ������������������������       �                     D@        .       7                     N@h�����?'             L@       /       0                   `l@      �?             @@       ������������������������       �                     5@        1       2                   �\@"pc�
�?	             &@        ������������������������       �                     �?        3       4                    �?ףp=
�?             $@       ������������������������       �                      @        5       6                    @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        ������������������������       �                     9@        ������������������������       �        +             Q@        ;       <                   @a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        >       o                   `a@ Р^D�?f            `d@       ?       P                    �?f<t=9%�?=             [@        @       O                    a@ZՏ�m|�?            �H@       A       B       
             �?��E�B��?            �G@        ������������������������       �                     @        C       L       	          033@�p ��?            �D@       D       E       	            �?�#-���?            �A@        ������������������������       �                     *@        F       G       	          ����?��2(&�?             6@        ������������������������       �                     �?        H       K                   �e@�����?             5@       I       J                   �`@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     �?        M       N                   �j@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        Q       \                   0l@TV����?             �M@        R       W       	          ����?l��
I��?             ;@       S       T                   `j@R���Q�?             4@        ������������������������       �                     &@        U       V                    �?�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        X       [                    �?����X�?             @       Y       Z                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ]       b                   �b@     ��?             @@        ^       a                   �`@���!pc�?             &@       _       `       	          ����?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        c       f       	          833�?����X�?             5@        d       e                   �^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        g       l                   �p@�r����?             .@       h       i                   pn@$�q-�?             *@       ������������������������       �                      @        j       k                    �F@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        m       n                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        p       �                    @lGts��?)            �K@       q       r       
             �?Hm_!'1�?$            �H@        ������������������������       �                     @        s       t                   0a@�����?             E@        ������������������������       �                     �?        u       ~                    �?��p\�?            �D@        v       }                    �?�r����?             .@       w       |                    �?      �?              @       x       {                    @M@؇���X�?             @        y       z                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               �       	          ����? ��WV�?             :@       ������������������������       �                     0@        �       �                    q@ףp=
�?             $@       ������������������������       �                      @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �j@�q�q�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                   pq@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    c@�#l��?�            �r@        �       �                    �?�	j*D�?             :@       �       �                    �?      �?             0@       �       �       	            �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �       	          033@<�N��?�            Pq@       �       �                    �?���"��?�            �p@       �       �                    �?`�c�г?�             o@        �       �                    �L@r�q��?'             K@       �       �                   @\@�ʈD��?            �E@        �       �                   �[@      �?	             (@       �       �                     E@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �       	          433�?�g�y��?             ?@       ������������������������       �                     8@        �       �                   �d@؇���X�?             @       ������������������������       �                     @        �       �                   0e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�eP*L��?             &@        �       �                    �?և���X�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �l@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @L@ �m�+�?t            @h@       ������������������������       �        b            �d@        �       �                   �_@ 7���B�?             ;@        �       �                    �L@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        �       �       	          433�?8�A�0��?             6@       �       �                   �r@ףp=
�?             $@       ������������������������       �                     @        �       �                   c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �E$�~V�?�����?�b�����?ZgND���?���[��?�_���@�?e�M6�d�?�M6�d��?�;�;�?'vb'vb�?              �?�;�;�?�؉�؉�?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?�������?      �?                      �?e�e��?��@��@�?�������?�������?C:o1��?��y�!�?br1���?g���Q��?w�qG��?⎸#��?���Q��?R���Q�?F]t�E�?/�袋.�?(�����?�k(���?              �?UUUUUU�?�������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?        9/���?������?      �?        UUUUUU�?UUUUUU�?              �?�$I�$I�?�m۶m��?      �?      �?              �?F]t�E�?/�袋.�?      �?        �������?�������?              �?      �?      �?              �?      �?                      �?              �?              �?      �?      �?              �?      �?        f5�8t�?�L����?����K�?������?9/����?�>4և��?AL� &W�?�l�w6��?              �?��+Q��?Q��+Q�?_�_�?�A�A�?              �?t�E]t�?��.���?      �?        �a�a�?=��<���?�������?ffffff�?              �?      �?              �?              �?      �?      �?                      �?      �?        E�pR���?u_[4�?Lh/����?h/�����?333333�?333333�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?                      �?      �?              �?      �?F]t�E�?t�E]t�?�q�q�?�q�q�?              �?      �?                      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?        �?�������?;�;��?�؉�؉�?              �?�������?�������?              �?      �?              �?      �?              �?      �?        �־a�?�<%�S��?9/���?Y�Cc�?              �?�a�a�?=��<���?      �?        ��+Q��?�]�ڕ��?�?�������?      �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?                      �?;�;��?O��N���?              �?�������?�������?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �I��A��?��be�F�?;�;��?vb'vb'�?      �?      �?�������?�������?      �?                      �?              �?              �?m�ǈ�?��� ù�?c��)F�?�\y@�ε?��Zk���?��RJ)��?�������?UUUUUU�?A_���?�}A_з?      �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?��{���?�B!��?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        t�E]t�?]t�E�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?:*����?���u?      �?        	�%����?h/�����?�������?UUUUUU�?              �?      �?              �?        /�袋.�?颋.���?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�A�'hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK˅�h��B�2         �                   �b@j8je3�?�           ��@              c       
             �?�+��8�?B           `@                                 �Y@�$���?�            �v@                      
             �?���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @               :                    �?�����H�?�            �u@              #       	          ����?($�pa�?�            q@        	                          �s@�����?E            �Z@       
                           �? i���t�?@            �X@                                  �?r�q��?)             N@                                 �p@L紂P�?"            �I@                     	          ����?H�V�e��?             A@       ������������������������       �                     8@                                  `_@�z�G��?             $@                                 �\@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             1@                                  �X@�q�q�?             "@        ������������������������       �                     �?                                  �]@      �?              @        ������������������������       �                     @                                  @_@�q�q�?             @        ������������������������       �                     �?                                  �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     C@               "                   ��@      �?              @               !                    ]@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        $       '                    �?��Q���?c            �d@        %       &                    f@ףp=
�?
             4@        ������������������������       �                      @        ������������������������       �        	             2@        (       /       
             �?@�E�x�?Y            `b@        )       .       	          ��� @HP�s��?             9@        *       -                   @\@"pc�
�?             &@        +       ,                    b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ,@        0       1                    �? ��7��?J            �^@       ������������������������       �        :             X@        2       3       	             @ ��WV�?             :@       ������������������������       �                     1@        4       9       	             @�����H�?             "@       5       8                    �?r�q��?             @       6       7                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ;       X                    �?����?4            �S@        <       S                    �?\�Uo��?             C@       =       >       
             �?      �?             <@        ������������������������       �                     @        ?       F                   @g@� �	��?             9@        @       E                   @b@�<ݚ�?             "@       A       D                    @K@      �?              @        B       C                    \@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        G       H                    �?      �?             0@        ������������������������       �                     @        I       J                    �?�q�q�?	             (@        ������������������������       �                     �?        K       L                   0b@���!pc�?             &@        ������������������������       �                     @        M       R                     P@���Q��?             @       N       Q                    `@      �?             @       O       P                   pn@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        T       W                    �?ףp=
�?             $@        U       V                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        Y       b                    �?ףp=
�?             D@       Z       [                    @M@؇���X�?             <@        ������������������������       �                     *@        \       a                    �?������?             .@       ]       `                     N@8�Z$���?	             *@        ^       _       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     (@        d                           �?T�iA�?a            �a@        e       n       	          ����?����"�?*             M@       f       m                     P@�����H�?             B@       g       h                     L@Pa�	�?            �@@       ������������������������       �                     <@        i       j       	          ����?z�G�z�?             @       ������������������������       �                     @        k       l                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       v                    �?"pc�
�?             6@        p       q       	          ����?���Q��?             @        ������������������������       �                      @        r       s       	          `ff�?�q�q�?             @        ������������������������       �                     �?        t       u                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        w       z                    �?�t����?             1@        x       y                   0a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        {       |                   �b@@4և���?
             ,@       ������������������������       �                     (@        }       ~                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @c@��1��?7            �T@        �       �                    �?�����H�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �_@���(-�?3            @R@        �       �                   �p@�����H�?             ;@       ������������������������       �                     5@        �       �                   Hq@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        "             G@        �       �       	             @���Bb�?�             m@       �       �       
             �?nғzw)�?�            �j@        �       �                    �?�;�vv��?*            @R@        �       �       	          ����?      �?             8@       ������������������������       �        	             &@        �       �                   �a@��
ц��?             *@       �       �                    �?���Q��?             $@       �       �                    �?�q�q�?             "@       �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �                   �r@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?f�Sc��?            �H@       �       �       	          ����?^����?            �E@       �       �                   `]@r�q��?             8@        ������������������������       �                      @        �       �                   `m@�C��2(�?             6@        ������������������������       �                     &@        �       �                   �m@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �G@D�n�3�?             3@        ������������������������       �                     @        �       �                   Pl@և���X�?             ,@        �       �                    �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�-x�j�?Z            `a@        �       �                    �L@�lg����?            �E@       �       �                    `@�������?             A@        �       �                   �c@���|���?             &@        ������������������������       �                     @        �       �                    �I@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �c@���}<S�?             7@        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             3@        �       �       	          ����?�<ݚ�?             "@       �       �                    �N@      �?              @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �t@p�qG�??             X@       ������������������������       �        :            �U@        �       �                   u@      �?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             4@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ���Y��?t�S��?��.�*��?����.�?"H��h��?����e��?F]t�E�?t�E]t�?              �?      �?        �q�q�?�q�q�?,�,��?~ڧ}ڧ�?5�x+��?��!5�x�?����X�?/�����?UUUUUU�?�������?�������?�������?ZZZZZZ�?iiiiii�?              �?ffffff�?333333�?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?      �?�m۶m��?�$I�$I�?              �?      �?                      �?\��l���?K��
�?�������?�������?      �?                      �?9/���?և���X�?{�G�z�?q=
ףp�?F]t�E�?/�袋.�?      �?      �?              �?      �?                      �?              �?;ڼOqɀ?��:ڼ�?              �?;�;��?O��N���?              �?�q�q�?�q�q�?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?��-��-�?H�4H�4�?6��P^C�?�5��P^�?      �?      �?      �?        )\���(�?�Q����?9��8���?�q�q�?      �?      �?      �?      �?              �?      �?              �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        t�E]t�?F]t�E�?              �?333333�?�������?      �?      �?      �?      �?              �?      �?              �?                      �?�������?�������?      �?      �?      �?                      �?              �?�������?�������?�$I�$I�?۶m۶m�?              �?�?wwwwww�?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?PuPu�?��+��+�?	�=����?�i��F�?�q�q�?�q�q�?|���?|���?      �?        �������?�������?      �?              �?      �?              �?      �?                      �?F]t�E�?/�袋.�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �?<<<<<<�?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?        �+Q���?,Q��+�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?��իW��?�P�B�
�?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?        ��{a�?����=�?:�&oe�?����!5�?�8�?����Ǐ�?      �?      �?              �?�؉�؉�?�;�;�?333333�?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?����>�?������?�qG��?w�qG��?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?        /�袋.�?F]t�E�?              �?      �?        l(�����?(������?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?              �?��\*�?ݘ��V�?}A_��?�}A_��?�������?�������?F]t�E�?]t�E]�?              �?�������?�������?      �?                      �?ӛ���7�?d!Y�B�?      �?      �?      �?                      �?      �?        �q�q�?9��8���?      �?      �?              �?      �?      �?      �?                      �?      �?        UUUUUU�?�������?      �?              �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK兔h��B@9         �       
             �?�^�P��?�           ��@                                  @G@r�g�?
           �z@                                  �n@     x�?'             P@              	                   �`@�K��&�?            �E@                                  pb@@4և���?
             ,@       ������������������������       �                     (@                                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        
                          �Q@д>��C�?             =@        ������������������������       �                      @                                   @�����H�?             ;@                                 `a@$�q-�?             :@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �? �q�q�?             8@        ������������������������       �                     &@                                   �C@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     5@               Y                    �?��a�2��?�            �v@               $       	          833�?��
n��?U            �a@                                   �?@4և���?             E@       ������������������������       �                     <@                                   �?d}h���?             ,@                                    P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                #                   `X@�C��2(�?	             &@       !       "                   `X@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        %       ,                   �g@D��ٝ�?:            @Y@        &       '                    �? 	��p�?             =@       ������������������������       �        
             *@        (       +       	             �?      �?             0@       )       *       
             �?"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        -       B                   �`@)O���?(             R@        .       A                     Q@�������?             >@       /       4                    @H@�>4և��?             <@        0       3                   �o@���Q��?             @        1       2       	          433�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        5       8                   `[@���}<S�?             7@        6       7                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        9       :                    �?���N8�?             5@        ������������������������       �                     @        ;       @                    �L@      �?             0@       <       =                   @q@      �?              @       ������������������������       �                     @        >       ?                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        C       H                    �M@X�Cc�?             E@        D       G                   p@      �?             0@       E       F                   @a@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        I       J       	          pff�?���B���?             :@        ������������������������       �                     �?        K       R                    _@�J�4�?             9@        L       Q                    �?և���X�?             @       M       P                   �\@      �?             @       N       O                    `P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        S       T                   pc@�X�<ݺ?             2@        ������������������������       �                     &@        U       V                   `a@؇���X�?             @        ������������������������       �                     �?        W       X                   �c@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       �                    �?��ҘR�?�             k@       [       x                   �_@ >�֕�?p            �e@       \       c                    �?�#-���?C            @Z@        ]       ^       
             �?�q�q�?             "@        ������������������������       �                      @        _       `                   �`@և���X�?             @        ������������������������       �                     �?        a       b                     L@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        d       u                   `_@      �?>             X@       e       f                   �i@`Ӹ����?:            �V@        ������������������������       �                     =@        g       t                   �a@��GEI_�?(            �N@       h       m       	          `ff�?��� ��?             ?@        i       l                    \@      �?	             (@        j       k                    `@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        n       o                    �?�}�+r��?             3@       ������������������������       �                     (@        p       q       	             @؇���X�?             @        ������������������������       �                     @        r       s                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@        v       w                   Pi@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        y       z                   `a@`����֜?-            �Q@        ������������������������       �                     @@        {       |                    @M@P�Lt�<�?             C@        ������������������������       �                     2@        }       �                    �M@P���Q�?             4@        ~                          `c@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        �       �                   �s@����X�?             E@       �       �                    �J@@�0�!��?             A@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?\-��p�?             =@       �       �                   �X@���y4F�?             3@        �       �                   0m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �M@      �?             0@        ������������������������       �                     @        �       �                   �`@�<ݚ�?	             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             $@        �       �                   xt@      �?              @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�s�$$��?�            `s@       �       �                    @L@���:�?�            pp@       �       �                    �?(;L]n�?�            @j@        �       �       	          033@�?�P�a�?&             N@       �       �                   @E@�j��b�?%            �M@        �       �                    �?      �?             @       �       �                   �X@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `\@,�+�C�?!            �K@        �       �                   �q@������?	             .@       �       �                   �l@d}h���?             ,@       �       �                    �?      �?              @        ������������������������       �                     �?        �       �                     I@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     D@        ������������������������       �                     �?        ������������������������       �        c            �b@        �       �                   �s@`��}3��?'            �J@       �       �                    @N@��+7��?"             G@        �       �                    �?�û��|�?             7@        ������������������������       �                     @        �       �                   @k@�\��N��?             3@       �       �                   �`@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �L@      �?              @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   Pn@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�LQ�1	�?             7@       ������������������������       �                     3@        �       �                   �_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �a@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   u@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �[@z�J��?            �G@        ������������������������       �                     @        �       �                    f@�>$�*��?            �D@       �       �                   �a@��+��?            �B@       �       �                    �?��}*_��?             ;@        �       �                   �^@�����H�?             "@        �       �       	          833�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             2@       �       �                   a@�q�q�?
             (@        �       �                   @a@���Q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   ht@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @b@r�q��?             @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �Z@ףp=
�?             $@        �       �                     L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�b��
     h�h)h,K ��h.��R�(KK�KK��hb�BP  ��1W-��?�<gTi��?�!5�x+�?����!5�?      �?     ��?��)kʚ�?���)k��?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?        a���{�?|a���?              �?�q�q�?�q�q�?�؉�؉�?;�;��?      �?      �?              �?      �?        �������?UUUUUU�?      �?        �؉�؉�?;�;��?              �?      �?                      �?              �?�q�q�?��8��8�?���G�>�?9 2ܫ`�?�$I�$I�?n۶m۶�?              �?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?]t�E�?�������?�������?      �?                      �?              �?z��~�X�?�7���S�?�{a���?������?              �?      �?      �?F]t�E�?/�袋.�?      �?                      �?              �?9��8���?��8��8�?�������?�������?�$I�$I�?�m۶m��?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?ӛ���7�?d!Y�B�?      �?      �?              �?      �?        ��y��y�?�a�a�?      �?              �?      �?      �?      �?      �?              �?      �?              �?      �?              �?                      �?�m۶m��?%I�$I��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        ى�؉��?��؉���?      �?        {�G�z�?�z�G��?۶m۶m�?�$I�$I�?      �?      �?      �?      �?              �?      �?              �?                      �?�q�q�?��8��8�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?      �?                      �?��g�3��?��y��?�A�A�?��+��+�?_�_�?�A�A�?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?l�l��??�>��?              �?;ڼOqɰ?�d����?�B!��?�{����?      �?      �?333333�?�������?              �?      �?                      �?(�����?�5��P�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�A�A�?�������?              �?(�����?���k(�?              �?�������?ffffff�?UUUUUU�?�������?      �?                      �?              �?�$I�$I�?�m۶m��?�������?ZZZZZZ�?�������?333333�?      �?                      �?�{a���?a����?(������?6��P^C�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?�q�q�?9��8���?              �?      �?                      �?      �?      �?      �?                      �?�����?�=���?����p�?H�x\�?�������?�?DDDDDD�?�����ݽ?�N��?��/���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�}��7��?��)A��?wwwwww�?�?I�$I�$�?۶m۶m�?      �?      �?              �?�m۶m��?�$I�$I�?      �?                      �?      �?                      �?      �?                      �?      �?        �琚`��?M0��>��?zӛ����?Y�B��?8��Moz�?��,d!�?      �?        y�5���?�5��P�?F]t�E�?t�E]t�?              �?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?      �?        ��Moz��?Y�B��?      �?              �?      �?      �?                      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        }g���Q�?AL� &W�?              �?�18���?�����?�S�n�?*�Y7�"�?B{	�%��?_B{	�%�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        �������?�������?      �?      �?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJJ��hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         �                    �?(��e��?�           ��@              7                    �J@$/2�l��?           P{@                      
             �?�LQ�1	�?l             d@                                  �?Hm_!'1�?D            �X@              
                   `m@�?�<��?1            @P@               	                   �f@ �q�q�?             8@                                  `U@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        	             *@                                   �?��r._�?!            �D@                                   �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @                                   @H@l��\��?             A@       ������������������������       �                     4@                                  `^@d}h���?             ,@        ������������������������       �                      @                      	             @�8��8��?
             (@       ������������������������       �                     "@                                   @J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �@@               0                    e@���N8�?(            �O@              %                    @F@�q�q�?             H@                                   �c@j���� �?             1@                                 pb@���!pc�?             &@                                    E@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        !       "                    �?�q�q�?             @        ������������������������       �                     �?        #       $                   �g@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        &       /                   �d@��� ��?             ?@       '       .                   �_@ףp=
�?             >@        (       +                    �?     ��?             0@        )       *                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ,       -       	          ����?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     �?        1       2                   �e@��S�ۿ?	             .@        ������������������������       �                     @        3       4                    �?      �?              @       ������������������������       �                     @        5       6                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        8       q       	             �?�A����?�            @q@        9       R       
             �?���y4F�?P            �`@       :       M                   `b@��� ��?9            @W@       ;       J                   pt@�����?2             U@       <       =                   �g@XI�~�?/            @S@       ������������������������       �                     C@        >       I                    �?�ݜ�?            �C@       ?       B                     L@���B���?             :@        @       A                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        C       D                   �[@�LQ�1	�?             7@        ������������������������       �                     �?        E       H                    �?�C��2(�?             6@        F       G                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     *@        K       L                     L@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        N       O       	            �?X�<ݚ�?             "@        ������������������������       �                     @        P       Q                    d@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        S       j                    �?���Q��?             D@       T       i                   `u@�q�q�?            �@@       U       d                    �?>���Rp�?             =@       V       Y                    �?ҳ�wY;�?	             1@        W       X                     N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       c                   d@�n_Y�K�?             *@       [       b       	             �?����X�?             @       \       a                    �?���Q��?             @       ]       ^                   �l@      �?             @        ������������������������       �                      @        _       `                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        e       f                    �N@�8��8��?             (@       ������������������������       �                     @        g       h                   �s@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        k       p       	             �?����X�?             @       l       o                    T@�q�q�?             @        m       n                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        r       �                    �?��K˱F�?S            �a@       s       x                   @^@@��j$޷?=            �Y@        t       u       	          `ff�?z�G�z�?             $@        ������������������������       �                     �?        v       w                   �]@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        y       ~                   �b@hl �&�?6             W@       z       }       	          ����? }�Я��?4            @V@        {       |                    c@�}�+r��?             3@       ������������������������       �        
             2@        ������������������������       �                     �?        ������������������������       �        )            �Q@               �                    @N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �D@        �       �                    �?:ɨ��?�            �r@        �       �                    `@�8��8N�?C             X@       �       �                    �K@ pƵHP�?#             J@       ������������������������       �                    �G@        �       �       
             �?z�G�z�?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @L@��2(&�?              F@       �       �                    �?(;L]n�?             >@       ������������������������       �                     ;@        �       �                    �J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    @O@X�Cc�?             ,@        �       �                   po@����X�?             @       �       �                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?��0��?�             i@        �       �       	          ���@��~l�?@            @V@       �       �                    �F@RB)��.�??            �U@        �       �                    @�q�q�?	             (@       �       �                    �C@      �?              @       �       �                   �r@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��A��?6            �R@        �       �                    �?X�Cc�?             ,@        �       �                    @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    `P@և���X�?             @       �       �       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   pk@�r����?*             N@       �       �                   @e@�IєX�?             A@       �       �                    �?�g�y��?             ?@        �       �                    �?$�q-�?             *@       ������������������������       �                     "@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �a@�θ�?             :@       ������������������������       �        	             *@        �       �                    �I@��
ц��?             *@        ������������������������       �                     @        �       �       	          ����?      �?              @       ������������������������       �                     @        �       �                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @������?G             \@       �       �       	            �?ܴD��?C            @Y@       ������������������������       �        :            @U@        �       �                    �?      �?	             0@       �       �                    �M@���!pc�?             &@       �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �U@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	             @�eP*L��?             &@       �       �                   pg@      �?              @        ������������������������       �                     @        �       �                    �J@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  M��+��?ڸ�j�?�t�	��?ۢ�=�{�?d!Y�B�?Nozӛ��?9/���?Y�Cc�? �����?�����?UUUUUU�?�������?F]t�E�?]t�E�?              �?      �?                      �?ە�]���?�ڕ�]��?�$I�$I�?۶m۶m�?      �?                      �?�������?------�?              �?۶m۶m�?I�$I�$�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�a�a�?��y��y�?�������?�������?ZZZZZZ�?�������?t�E]t�?F]t�E�?333333�?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?        �{����?�B!��?�������?�������?      �?      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?�?      �?              �?      �?      �?              �?      �?      �?                      �?�Mozӛ�?C���,�?(������?6��P^C�?�B!��?�{����?�a�a�?=��<���?V~B����?5�wL��?              �?�i�i�?\��[���?ى�؉��?��؉���?UUUUUU�?UUUUUU�?              �?      �?        Y�B��?��Moz��?      �?        F]t�E�?]t�E�?�������?333333�?              �?      �?                      �?              �?۶m۶m�?�$I�$I�?              �?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?GX�i���?�i��F�?�������?�������?      �?      �?      �?                      �?ى�؉��?;�;��?�m۶m��?�$I�$I�?333333�?�������?      �?      �?      �?              �?      �?      �?                      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �L[���?0K����?�?nnnnnn�?�������?�������?      �?        �q�q�?�q�q�?      �?                      �?Y�B��?ozӛ���?p�\��?�я~���?(�����?�5��P�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?N6�d�M�?e�M6�d�?�������?�������?'vb'vb�?;�;��?      �?        �������?�������?      �?      �?      �?                      �?      �?        ��.���?t�E]t�?�������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?%I�$I��?�m۶m��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        b�V�;��?<�RG�m�?��x�3�?�9�as�?���)k��?S֔5eM�?�������?�������?      �?      �?      �?      �?              �?      �?              �?                      �?�g�`�|�?��g�`�?�m۶m��?%I�$I��?�$I�$I�?۶m۶m�?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?        �?�������?�?�?�B!��?��{���?;�;��?�؉�؉�?              �?      �?      �?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?ى�؉��?              �?�؉�؉�?�;�;�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        n۶m۶�?I�$I�$�?�(0���?z��~�X�?      �?              �?      �?t�E]t�?F]t�E�?�q�q�?�q�q�?              �?      �?              �?        333333�?�������?              �?      �?        t�E]t�?]t�E�?      �?      �?      �?        333333�?�������?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�U�uhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�.         h                    �?8}�ý�?�           ��@              E       
             �?|�e4@@�?           �{@                                   �G@r%����?s            �f@               	                    �?h+�v:�?             A@                                   �D@r�q��?             (@       ������������������������       �                     "@                                   @F@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        
                          0o@��2(&�?             6@       ������������������������       �                     2@                                   �?      �?             @        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                      	          ����?B`�I��?\            `b@                                  �b@���N8�?             E@       ������������������������       �                    �A@                                  `a@����X�?             @       ������������������������       �                     @        ������������������������       �                      @                       	          ����?^������?A            @Z@                                  0c@���N8�?             5@       ������������������������       �                     (@                                  @a@X�<ݚ�?             "@                                   �J@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �N@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        !       D                    @R@���N8�?4             U@       "       3                   �b@��P���?3            �T@       #       ,                   0b@�8��8��?#             N@       $       )                   xr@ �q�q�?             H@       %       (                   �^@����?�?            �F@        &       '                    �P@      �?	             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     =@        *       +                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        -       2                   �`@      �?             (@       .       1                   @q@      �?              @       /       0       	          033�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        4       A                   `d@8�A�0��?             6@       5       <       	             @      �?             0@       6       7       	          033�?�8��8��?             (@       ������������������������       �                     @        8       ;                    �K@r�q��?             @       9       :       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        =       >                   �c@      �?             @        ������������������������       �                      @        ?       @                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        B       C                    b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        F       g       	          `ff@8�����?�            �p@       G       Z                    �?�Wz��?�            0p@        H       W       	          ����?���N8�?&            �O@       I       T                    b@"pc�
�?             �K@       J       M                   @E@L紂P�?            �I@        K       L       	          ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        N       S                    ]@���}<S�?             G@        O       P                   �b@����X�?             ,@       ������������������������       �                     "@        Q       R                   �c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @@        U       V                    �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        X       Y       	          ����?      �?              @        ������������������������       �                     @        ������������������������       �                     @        [       f                     R@ %$��ݞ?u            �h@       \       ]                     L@@�[0)ʔ?t            `h@       ������������������������       �        [             c@        ^       e       	          ����?���N8�?             E@       _       `                   �b@�8��8��?             8@        ������������������������       �                     *@        a       b                    �L@"pc�
�?             &@        ������������������������       �                     �?        c       d                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        
             2@        ������������������������       �                     �?        ������������������������       �                     @        i       �       	          ����?x�>}��?�            �q@        j       s                    l@�q����?(            �J@       k       r                    �L@`Jj��?             ?@        l       q                    �?r�q��?             (@       m       p                    �K@z�G�z�?             $@       n       o                   Pj@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        t       u                   �l@���|���?             6@        ������������������������       �                     @        v       y                    �?X�<ݚ�?             2@        w       x                   pb@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        z       �                    b@�q�q�?	             (@       {       �                    @L@X�<ݚ�?             "@       |       �       	          ����?�q�q�?             @       }       �                    �H@z�G�z�?             @       ~                           ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �R@$�q-�?�            @m@       �       �                    Z@��ۆ�P�?�             m@        �       �                   �Y@      �?              @       �       �                    �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?Х-��ٹ?�             l@       �       �                    @E@ 7���B�?e            @d@        �       �       
             �?8�Z$���?
             *@        ������������������������       �                     �?        �       �                    �D@r�q��?	             (@       �       �                    �C@�C��2(�?             &@       ������������������������       �                      @        �       �                   �i@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �? �ޫ��?[            �b@       �       �                   `a@�����?R             a@        ������������������������       �        (            �O@        �       �       	             @���(-�?*            @R@       �       �                   �b@�1�`jg�?!            �K@       �       �                   �b@���J��?            �I@       ������������������������       �                     ;@        �       �                    �? �q�q�?             8@       ������������������������       �                     7@        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             2@        �       �                    �?$�q-�?	             *@        �       �                   �`@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    c@�����?&            �O@       �       �                    �?�X�<ݺ?              K@       �       �                   0p@���.�6�?             G@       �       �                   �X@      �?             @@        ������������������������       �                     �?        ������������������������       �                     ?@        �       �                   �_@؇���X�?             ,@        �       �                    @J@���Q��?             @        ������������������������       �                      @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        �       �                     L@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  a[ӿc�?PR Np�?ExR��y�?w[��?������?2������?�������?xxxxxx�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?��.���?t�E]t�?      �?              �?      �?              �?      �?      �?      �?                      �?#��Q��?�(W��?�a�a�?��y��y�?              �?�$I�$I�?�m۶m��?              �?      �?        _�_��?uPuP�?�a�a�?��y��y�?      �?        �q�q�?r�q��?      �?      �?      �?                      �?�������?�������?              �?      �?        ��y��y�?�a�a�?�����?������?UUUUUU�?UUUUUU�?UUUUUU�?�������?l�l��?��I��I�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?      �?      �?              �?      �?                      �?              �?颋.���?/�袋.�?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?      �?      �?                      �?UUUUUU�?�������?              �?      �?              �?        �τ?��?���f�?k�����?���ʱ?�a�a�?��y��y�?/�袋.�?F]t�E�?�������?�������?�������?333333�?      �?                      �?ӛ���7�?d!Y�B�?�m۶m��?�$I�$I�?      �?        �������?�������?              �?      �?              �?              �?      �?      �?                      �?      �?      �?              �?      �?        ������?և���X�?�������?PP�?      �?        ��y��y�?�a�a�?UUUUUU�?UUUUUU�?      �?        /�袋.�?F]t�E�?              �?�������?�������?              �?      �?              �?                      �?              �?�B���S�?����5�?�x+�R�?�Cj��V�?�B!��?���{��?UUUUUU�?�������?�������?�������?�q�q�?�q�q�?              �?      �?              �?                      �?              �?]t�E]�?F]t�E�?      �?        r�q��?�q�q�?�������?UUUUUU�?              �?      �?        �������?�������?r�q��?�q�q�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?              �?                      �?;�;��?�؉�؉�?�l�����?gR��L��?      �?      �?�������?333333�?              �?      �?              �?        O贁N�?K~��K�?h/�����?	�%����?;�;��?;�;��?              �?UUUUUU�?�������?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �3�=l}�?d.�$�?�������?KKKKKK�?              �?�P�B�
�?��իW��?�־a�?A��)A�?�?______�?              �?UUUUUU�?�������?              �?      �?              �?      �?      �?                      �?              �?;�;��?�؉�؉�?UUUUUU�?�������?      �?                      �?              �?�a�a�?=��<���?�q�q�?��8��8�?Y�B��?���7���?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW��]hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�/         B                   �_@6�L����?�           ��@               !                    �?����k�?�            Pp@                                   �?k��9�?;            �V@                                 �^@Nd^����?)            �N@                                 �\@�q�q�?$            �I@                                  U@�'�=z��?            �@@        ������������������������       �                     @                                   �?�f7�z�?             =@       	                          �Y@և���X�?             5@        
                           @L@      �?              @       ������������������������       �                     @                                   @      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                  @i@�	j*D�?
             *@        ������������������������       �                     @                      	             �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                  @^@�X�<ݺ?             2@       ������������������������       �        	             .@                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                   �?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @                                  �n@ 	��p�?             =@       ������������������������       �                     :@                       	          033�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        "       =       
             �?�E}�<>�?k            `e@       #       :                   `f@ �&�eZ�?b             c@       $       9                   ``@x�C����?`            �b@        %       &       
             �?�8��8��?(             N@        ������������������������       �                     ,@        '       6       	          033@�q��/��?              G@       (       1                    �?���N8�?             E@       )       *                    �?�?�|�?            �B@        ������������������������       �                     $@        +       0                   �Z@ 7���B�?             ;@        ,       -                   �m@�8��8��?             (@       ������������������������       �                      @        .       /       	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        2       5                   �X@z�G�z�?             @        3       4                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        7       8                   �r@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        8             V@        ;       <                   �^@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        >       ?                   �[@b�2�tk�?	             2@        ������������������������       �                     @        @       A       	          ����?�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        C       �                    �?>^�3���?(           �}@       D       �       	          ���@��%�}�?�            �w@       E       ~       
             �?�+�Y��?�            0u@        F       e                   �b@+Y���?K            @\@       G       T                    �?:ɨ��?-            �P@        H       M                   Pa@��S���?             >@        I       J                    �?8�Z$���?             *@        ������������������������       �                     �?        K       L                    @D@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        N       O                   �\@@�0�!��?
             1@        ������������������������       �                     @        P       Q                    l@�z�G��?             $@        ������������������������       �                     @        R       S                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        U       Z                    �E@r�q��?             B@        V       Y                    `@      �?             @       W       X       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        [       d       	          ����?      �?             @@       \       c                    @r�q��?             8@       ]       ^                   �\@�LQ�1	�?             7@        ������������������������       �                      @        _       `                    f@���N8�?             5@       ������������������������       �                     2@        a       b                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        f       i                    �C@p�v>��?            �G@        g       h                   s@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        j       s                    @L@��P���?            �D@       k       r                    �? �Cc}�?             <@       l       q                   �b@�>����?             ;@       m       p                    �? ��WV�?             :@        n       o                    �G@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     �?        ������������������������       �                     �?        t       {                    �?��
ц��?             *@       u       v                    �?      �?             $@        ������������������������       �                     @        w       x                     @r�q��?             @        ������������������������       �                     @        y       z                   p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        |       }                   0p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               �                    �? (��?�            @l@        �       �                    ]@��s����?(            �O@        �       �                    �?�IєX�?	             1@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        �       �                    �?�5��
J�?             G@       �       �                    �?l��\��?             A@        �       �                    �G@      �?              @        ������������������������       �                      @        �       �                   �b@r�q��?             @       ������������������������       �                     @        �       �                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        �       �                   a@�q�q�?	             (@        ������������������������       �                      @        �       �                     M@z�G�z�?             $@       �       �                   @d@      �?              @       �       �       	             �?؇���X�?             @       �       �                   �b@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    d@�dJ�Ҙ?c            `d@       ������������������������       �        4             X@        �       �                     L@0�,���?/            �P@       ������������������������       �        (            �M@        �       �                   �m@      �?              @        �       �                    e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �j@�?�|�?            �B@        �       �                    @H@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     =@        �       �       
             �?�E���?<            @X@       �       �                    �?(��+�?'            �N@       ������������������������       �                     D@        �       �       	          ����?�ՙ/�?             5@        ������������������������       �                     @        �       �                     K@      �?
             0@        ������������������������       �                     @        �       �       	          ����?�n_Y�K�?             *@        ������������������������       �                     @        �       �       	          ����?�����H�?             "@        ������������������������       �                     @        �       �       	          ��� @�q�q�?             @       �       �                    p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          033�?�<ݚ�?             B@       �       �                   �r@XB���?             =@       ������������������������       �                     ;@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  6�;����?e���?��B�}��?_S����?[�[��?�'}�'}�?�u�y���?���:�?UUUUUU�?UUUUUU�?|��|�?|���?              �?O#,�4��?a���{�?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?              �?      �?        ;�;��?vb'vb'�?              �?�q�q�?r�q��?      �?                      �?      �?        ��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?�{a���?������?              �?UUUUUU�?UUUUUU�?      �?                      �?XOa=���?�SXOa�?�l�l�?�3��3��?���L�?�n0E>��?UUUUUU�?UUUUUU�?              �?��Mozӻ?�B����?�a�a�?��y��y�?к����?*�Y7�"�?              �?h/�����?	�%����?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?�������?�������?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?              �?�������?333333�?              �?      �?        9��8���?�8��8��?              �?�������?�������?      �?                      �?3ru�hn�?�.#�?��F}g��?br1��?j<����?Y�����?H���?��	���?e�M6�d�?N6�d�M�?�������?�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?ZZZZZZ�?              �?333333�?ffffff�?              �?      �?      �?      �?                      �?UUUUUU�?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?UUUUUU�?�������?Y�B��?��Moz��?      �?        �a�a�?��y��y�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?ڨ�l�w�?L� &W�?UUUUUU�?�������?              �?      �?        ������?�����?%I�$I��?۶m۶m�?�Kh/��?h/�����?O��N���?;�;��?      �?      �?      �?                      �?      �?                      �?              �?�;�;�?�؉�؉�?      �?      �?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        H���?x�!���?z��y���?�a�a�?�?�?      �?      �?      �?                      �?      �?        �,d!Y�?�Mozӛ�?------�?�������?      �?      �?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?�������?      �?                      �?              �?      �?                      �?w��|��?)��I� �?      �?        Ez�rv�?g��1��?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        к����?*�Y7�"�?      �?      �?      �?                      �?              �?W?���?tT����?;ڼOq��?q�����?              �?�a�a�?�<��<��?              �?      �?      �?      �?        ى�؉��?;�;��?      �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?9��8���?�q�q�?GX�i���?�{a���?      �?              �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJt�mUhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKǅ�h��B�1         V       	             �?n3�ԉ[�?�           ��@               7                    �?d%@�"�?�            �u@                                  �[@DX�\��?_            �a@               	                   `V@��G���?            �B@                                 �Z@ 7���B�?             ;@       ������������������������       �                     5@                                   [@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        
                          �Z@���Q��?	             $@                                   �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  0k@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  pi@��
P��?F            @Z@                                  0g@      �?             D@                                  �?�n_Y�K�?             :@                                 @E@X�<ݚ�?             2@                                  �Z@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   _@"pc�
�?             &@        ������������������������       �                     �?                                   �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@               2       	          833�?�7�֥��?,            @P@               !       
             �?<|ۤ$�?$            �K@        ������������������������       �                     &@        "       '                    �I@���!pc�?             F@       #       &                    �?�����?             5@       $       %                     B@�����H�?             2@        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     @        (       -                   �c@\X��t�?             7@        )       *       	          ����?�8��8��?             (@       ������������������������       �                     $@        +       ,                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        .       /                   Pd@"pc�
�?             &@       ������������������������       �                      @        0       1                   �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        3       6                   �_@ףp=
�?             $@        4       5                    r@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        8       G       
             �?~�4��m�?�             j@        9       >                    @H@l`N���?            �J@        :       ;                    @C@z�G�z�?	             .@        ������������������������       �                      @        <       =                    �?$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ?       F                    �O@�d�����?             C@       @       A       
             �?z�G�z�?            �A@        ������������������������       �                     @        B       E                   �_@XB���?             =@        C       D       	          ����?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     @        H       I                    @L@�7��?i            �c@       ������������������������       �        X             `@        J       S                   �s@����X�?             <@       K       P                    c@��2(&�?             6@       L       M                   �a@�}�+r��?             3@        ������������������������       �                     (@        N       O                   0b@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        Q       R       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        T       U                    `@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        W       �                   a@��[̖x�?�            �w@       X       �       
             �?�Ӆ�0�?�            `m@       Y       r                   P`@��a�n`�?}             k@        Z       m                   8r@������?1            �V@       [       `                   �i@�Zl�i��?,            @T@        \       ]                    @O@`���i��?             F@       ������������������������       �                     C@        ^       _                    `@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        a       j       	          033@��G���?            �B@       b       e                    �?      �?             @@        c       d                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        f       i                   `X@ ��WV�?             :@        g       h                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        k       l                   @^@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        n       o                    �?�z�G��?             $@        ������������������������       �                     �?        p       q                    ]@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        s       v                    �D@���N8�?L            �_@        t       u       	             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        w       �                    @ ;=֦��?J            �^@       x       }                    �R@ �.�?Ƞ?H             ^@       y       |                    �?�6H�Z�?F            @]@        z       {                    �?�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �        =            @Z@        ~              
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �u@�E��ӭ�?             2@       �       �                    �?������?             1@       �       �                    �?�8��8��?
             (@        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                   �b@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?����-�?[            �b@        �       �       
             �?�G�V�e�?(             Q@        ������������������������       �                     *@        �       �                    �?�2����?!            �K@       �       �                   �\@�������?             A@        ������������������������       �                     @        �       �                    @F@r�q��?             >@        ������������������������       �                     �?        �       �                     M@\-��p�?             =@        ������������������������       �                     ,@        �       �                    �M@������?             .@        ������������������������       �                     �?        �       �                    �?d}h���?
             ,@        �       �       	          033	@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     5@        �       �                    �L@��Q��?3             T@       �       �                    �?�+e�X�?             I@        ������������������������       �                     "@        �       �                   �d@������?            �D@        ������������������������       �                     @        �       �       	             @���@��?            �B@       �       �                   �c@��hJ,�?             A@       �       �       
             �?     ��?             @@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    a@��S�ۿ?             >@       �       �                    �? 7���B�?             ;@        ������������������������       �                     (@        �       �       	          ����?��S�ۿ?	             .@        ������������������������       �                     @        �       �                    �?      �?              @       ������������������������       �                     @        �       �                   m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��S���?             >@        ������������������������       �                     @        �       �       
             �?�5��?             ;@       �       �                   o@      �?             2@       �       �                    �N@      �?             (@       �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�<ݚ�?             "@        ������������������������       �                      @        �       �                   �m@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  ����Gw�?��\D�?�LɔL��?�fm�fm�?�D+l$�?�]�����?v�)�Y7�?#�u�)��?h/�����?	�%����?              �?UUUUUU�?�������?      �?                      �?333333�?�������?�������?�������?      �?                      �?�������?333333�?              �?      �?        _�_��?PuPu�?      �?      �?ى�؉��?;�;��?r�q��?�q�q�?�$I�$I�?۶m۶m�?      �?                      �?/�袋.�?F]t�E�?              �?�������?�������?      �?                      �?              �?              �?�B/�B/�?z�z��?��)A��?��7�}��?              �?F]t�E�?t�E]t�?=��<���?�a�a�?�q�q�?�q�q�?              �?      �?              �?        !Y�B�?��Moz��?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?              �?      �?              �?        0��jY�?A۽U���?
�[���?�R���?�������?�������?              �?�؉�؉�?;�;��?      �?                      �?y�5���?Cy�5��?�������?�������?      �?        �{a���?GX�i���?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?        ��[��[�?�A�A�?      �?        �m۶m��?�$I�$I�?��.���?t�E]t�?�5��P�?(�����?      �?        ۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?      �?                      �?� �Ab�?տ�o'��?����R�?����u�?�c�1Ƹ?�s�9��?�Q�Q�?�������?�����H�?�"e����?F]t�E�?F]t�E�?              �?UUUUUU�?�������?      �?                      �?v�)�Y7�?#�u�)��?      �?      �?      �?      �?      �?                      �?;�;��?O��N���?      �?      �?              �?      �?                      �?333333�?�������?      �?                      �?ffffff�?333333�?              �?9��8���?�q�q�?              �?      �?        �a�a�?��y��y�?      �?      �?      �?                      �?XG��).�?�%C��6�?�?wwwwww�?���?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?r�q��?�q�q�?�?xxxxxx�?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?              �?      �?              �?        ��g�`�?��L���?�������?�������?              �?� O	��?��7�}��?�������?�������?      �?        UUUUUU�?�������?      �?        �{a���?a����?              �?�?wwwwww�?      �?        ۶m۶m�?I�$I�$�?      �?      �?      �?                      �?              �?              �?�������?ffffff�?R���Q�?���Q��?      �?        �v%jW��?��+Q��?              �?L�Ϻ��?к����?KKKKKK�?�������?      �?      �?      �?      �?              �?      �?        �������?�?	�%����?h/�����?      �?        �������?�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�?      �?        /�����?h/�����?      �?      �?      �?      �?�������?333333�?              �?      �?              �?                      �?�q�q�?9��8���?              �?�$I�$I�?�m۶m��?              �?      �?        �t�bub�G     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJc��hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         .                   �c@4�5����?�           ��@                      
             �?8�Z$���?e            �c@                                  �?4Qi0���?P            �^@                                   �?���B���?"             J@                                  �^@�n_Y�K�?             :@                                  �V@�n_Y�K�?             *@        ������������������������       �                     @               	                    �?z�G�z�?             $@        ������������������������       �                     @        
                           �M@      �?             @        ������������������������       �                      @        ������������������������       �                      @                      	          @33�?8�Z$���?             *@       ������������������������       �                     @                                  �d@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     :@                                  �e@ ��PUp�?.            �Q@       ������������������������       �        ,            @Q@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               -                    �?����e��?            �@@              &                    �?r�q��?             8@              !                    �?     ��?
             0@                                  @_@r�q��?             (@                                 `Y@�q�q�?             @        ������������������������       �                     �?                      	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        "       #                   �]@      �?             @        ������������������������       �                      @        $       %                    _@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        '       ,                   a@      �?              @       (       +                    �?      �?             @       )       *       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        /       j                   �`@�A�I���?k           �@        0       ;                   �h@.�Ȍ��?�            �l@        1       8                    �?���Q��?             >@       2       7                   @_@b�2�tk�?             2@       3       6       	             �?�8��8��?             (@        4       5                    �I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        9       :                     O@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        <       W       	          ����?�Tu�j��?x            �h@        =       B                    �?�o;����?3            �S@        >       ?                    �J@ףp=
�?             4@       ������������������������       �                     ,@        @       A                   `]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        C       P       
             �?TV����?&            �M@       D       E       
             �?R���Q�?             D@        ������������������������       �                      @        F       G       	          ����?>A�F<�?             C@       ������������������������       �                     2@        H       I                    �?��Q��?             4@        ������������������������       �                     @        J       K                    �O@@4և���?	             ,@       ������������������������       �                     $@        L       O                   �p@      �?             @       M       N                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        Q       V                    �O@�KM�]�?             3@       R       U                    �?�X�<ݺ?
             2@        S       T                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     �?        X       c                   �\@H��ԛ�?E            �]@        Y       ^                   �j@dP-���?             �G@        Z       ]                   ``@      �?              @        [       \                    @L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        _       b       
             �? ���J��?            �C@        `       a                   �r@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     A@        d       e                    @L@�k~X��?%             R@       ������������������������       �                     E@        f       i                    �L@(;L]n�?             >@        g       h       	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@        k       �       
             �?4��P8O�?�            �u@        l       s                   �a@.}Z*�?Z            �a@        m       n                    �?(;L]n�?             >@       ������������������������       �                     6@        o       r                    ^@      �?              @        p       q                   �n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       �       	          `ff@�Cc}��?F             \@       u       �                    �?h0�����?>            @Y@        v       �                    �?4�2%ޑ�?            �A@       w       x                     B@     ��?             @@        ������������������������       �                     �?        y       |                    �?��� ��?             ?@        z       {                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        }       �                   @^@ �q�q�?             8@        ~                           �K@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             1@        ������������������������       �                     @        �       �                    �?���e��?(            �P@       �       �       
             �?�G��l��?             E@        ������������������������       �                     @        �       �                   �[@b�2�tk�?             B@        ������������������������       �                     @        �       �                   xr@4���C�?            �@@       �       �                   0o@��X��?             <@       �       �                    �?���Q��?             .@       �       �                   �j@�	j*D�?
             *@        �       �                   @b@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �l@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     @        �       �                   �a@�q�q�?             8@        ������������������������       �                     @        �       �                    �?�d�����?
             3@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �H@�C��2(�?             &@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?4��?�?�             j@        �       �                   �b@     ��?'             P@        �       �                   `j@XB���?             =@        �       �                   `a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                    @I@�xGZ���?            �A@        �       �                    �?      �?
             0@        �       �                   �c@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                     G@ףp=
�?             $@       ������������������������       �                     @        �       �                    d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?p�ݯ��?             3@       �       �                   �c@��
ц��?	             *@        ������������������������       �                     @        �       �                   `a@�q�q�?             "@       �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                   �`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �t@@��8��?_             b@       �       �       	          ����?`����֜?[            �a@       �       �                    �? ��7��?O            �^@        �       �                     L@ �q�q�?             8@       ������������������������       �        
             4@        �       �                   `b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        B            �X@        �       �                    �?�X�<ݺ?             2@       ������������������������       �                     (@        �       �                    j@r�q��?             @        �       �                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?      �?             @        �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp   Np	�?���Gw{�?;�;��?;�;��?�On��?#6�a#�?ى�؉��?��؉���?ى�؉��?;�;��?;�;��?ى�؉��?              �?�������?�������?      �?              �?      �?              �?      �?        ;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?��V،?��ۥ���?              �?      �?      �?              �?      �?        6�d�M6�?e�M6�d�?UUUUUU�?UUUUUU�?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?߄*�u�?B��_��?�,�����?��,����?333333�?�������?9��8���?�8��8��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�~�@��?�R�֯�?�#{���?��	�Z�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        u_[4�?E�pR���?�������?�������?      �?        Cy�5��?������?              �?ffffff�?�������?      �?        �$I�$I�?n۶m۶�?              �?      �?      �?      �?      �?      �?                      �?              �?�k(���?(�����?��8��8�?�q�q�?      �?      �?      �?                      �?      �?                      �?:�:��?_̧^̧�?W�+�ɵ?�����F�?      �?      �?      �?      �?              �?      �?                      �?�A�A�?��-��-�?�������?�������?              �?      �?                      �?�q�q�?�8��8��?              �?�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?iȹ�. �?-o�`���?�
��V�?�z2~���?�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?�m۶m��?Q`ҩy�?�]?[��?�������?�A�A�?      �?      �?              �?�{����?�B!��?�$I�$I�?۶m۶m�?      �?                      �?�������?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?      �?                      �?>���>�?�>���?��y��y�?1�0��?      �?        9��8���?�8��8��?              �?'�l��&�?m��&�l�?%I�$I��?n۶m۶�?333333�?�������?vb'vb'�?;�;��?�������?333333�?      �?                      �?      �?      �?      �?              �?      �?      �?              �?      �?      �?                      �?              �?              �?      �?        �������?UUUUUU�?              �?y�5���?Cy�5��?      �?      �?              �?      �?        F]t�E�?]t�E]�?              �?      �?        F]t�E�?]t�E�?      �?      �?      �?                      �?              �?�N��N��?ى�؉��?     ��?      �?GX�i���?�{a���?      �?      �?              �?      �?              �?        �_�_�?�A�A�?      �?      �?      �?      �?              �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        Cy�5��?^Cy�5�?�;�;�?�؉�؉�?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?              �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?�������?�A�A�?��:ڼ�?;ڼOqɀ?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?        ��8��8�?�q�q�?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg�$hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKh��B�;         �                    �?6������?�           ��@              M       
             �?�)�@��?            z@                                  �`@���Q��?]             b@                                   �Q@�C��2(�?             F@                                  �?Du9iH��?            �E@                     
             �?(;L]n�?             >@        ������������������������       �                     @                                  �^@ �q�q�?             8@        	       
                   �Y@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             .@                                   �?8�Z$���?             *@                      	          `ff�?�q�q�?             @        ������������������������       �                     �?                                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  c@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?               (                    �?:�o���??            @Y@                                   �?*O���?             B@                                   �?      �?             $@                                 �a@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                    L@�	j*D�?             :@        ������������������������       �        	             $@                %                    �?      �?
             0@       !       $       	          `ff�?      �?             (@       "       #                   �\@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        &       '       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        )       *                    �A@�7�֥��?&            @P@        ������������������������       �                     @        +       ,                   `X@�BE����?%             O@        ������������������������       �                     @        -       2                    �G@��h!��?#            �L@        .       /                   0c@$�q-�?
             *@        ������������������������       �                     @        0       1                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        3       6                    �I@�X���?             F@        4       5                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        7       8       	          ����?�<ݚ�?             B@        ������������������������       �                     �?        9       F                   @c@z�G�z�?            �A@       :       ;                    �?      �?             8@        ������������������������       �                     $@        <       =                   @_@d}h���?	             ,@        ������������������������       �                     @        >       E                    @�z�G��?             $@       ?       B                    �?�<ݚ�?             "@       @       A                   @q@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        C       D                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        G       L                   @b@���|���?             &@       H       I                   d@�q�q�?             @        ������������������������       �                     @        J       K                   �o@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        N       _                    c@<Sw�[��?�            q@        O       P                     F@�	j*D�?             :@        ������������������������       �                     @        Q       V                    `@�ՙ/�?             5@        R       U                   �R@"pc�
�?             &@       S       T                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        W       \                    �L@���Q��?             $@       X       Y                    �?z�G�z�?             @        ������������������������       �                     @        Z       [                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                   �`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        `       o                    �?$�q-�?�            �n@        a       l                    �?�d�����?             C@       b       c                   �b@�LQ�1	�?             7@        ������������������������       �                     @        d       k                   Pe@      �?             0@       e       j                   ps@z�G�z�?             $@       f       g                    @H@�q�q�?             @        ������������������������       �                     @        h       i                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        m       n                   �e@�r����?
             .@       ������������������������       �        	             *@        ������������������������       �                      @        p       �                   �t@@�S�1�?}             j@       q       |                     L@�]��?z            �i@       r       s                    �?�B:�g�?e            �e@        ������������������������       �        &             M@        t       {                    �?@m���??             ]@       u       z                    ]@@��!�Q�?8            @Z@        v       y       	          ����?@4և���?             ,@       w       x                     I@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        0            �V@        ������������������������       �                     &@        }       �                    �M@     ��?             @@        ~                          �g@      �?              @        ������������������������       �                     �?        �       �       	          ����?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             8@        ������������������������       �                     $@        �       �                    �?d}h���?             ,@       �       �                    �N@�C��2(�?             &@        �       �                    @N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   (u@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �Y@(e����?�            �s@        ������������������������       �                     @        �       �                   i@8��#}N�?�            �s@        �       �                    �?�?�|�?B            �[@       ������������������������       �        0            @T@        �       �                   �e@ףp=
�?             >@       �       �       
             �? 	��p�?             =@       ������������������������       �                     3@        �       �                   �]@z�G�z�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@       �       �                   `b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �b@"����U�?�            @i@       �       �                    �?(��+�?u            �f@       �       �                    �?��a�n`�?a            `c@       �       �                   �a@؞�z�̼?F            @]@       �       �                    �?p=
ףp�?1             T@        ������������������������       �                     0@        �       �       	          ����?     ��?&             P@        �       �       	          ����?     ��?
             0@        �       �                    @G@      �?              @        ������������������������       �                     @        �       �                   �[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @K@      �?              @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   `_@ �q�q�?             H@        ������������������������       �                     6@        �       �                   `]@$�q-�?             :@        �       �                   �`@�q�q�?             @       �       �                    �K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     4@        ������������������������       �                    �B@        �       �                   (r@���y4F�?             C@       �       �                    m@ �Cc}�?             <@        ������������������������       �                     &@        �       �                   �`@@�0�!��?             1@       �       �       	             @�r����?
             .@       ������������������������       �                      @        �       �                    �?����X�?             @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             $@       �       �                   @^@����X�?             @       �       �       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          hff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��X��?             <@        ������������������������       �                     @        �       �       
             �?�㙢�c�?             7@       �       �                    �?��2(&�?             6@        �       �                    @      �?             @       �       �                   Pm@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����?�X�<ݺ?             2@        �       �       	             �?      �?             @        ������������������������       �                      @        �       �                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     �?        �       �                    �?D�n�3�?             3@       �       �                   �j@ҳ�wY;�?             1@        ������������������������       �                     @        �       �                    `@d}h���?             ,@        �       �                    �?և���X�?             @        ������������������������       �                      @        �       �                   �o@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��X�5�?��S�$e�?L"�Zց�?h��JS��?�������?333333�?F]t�E�?]t�E�?w�qGܱ?qG�w��?�?�������?              �?UUUUUU�?�������?�q�q�?�q�q�?      �?                      �?              �?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?�������?              �?      �?              �?        �g����?)0��<��?�q�q�?�q�q�?      �?      �?      �?      �?      �?                      �?              �?;�;��?vb'vb'�?              �?      �?      �?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?      �?      �?                      �?�B/�B/�?z�z��?              �?)��RJ)�?���Zk��?              �?Hp�}�?p�}��?�؉�؉�?;�;��?      �?        �������?UUUUUU�?      �?                      �?]t�E�?�E]t��?      �?      �?      �?                      �?9��8���?�q�q�?              �?�������?�������?      �?      �?      �?        I�$I�$�?۶m۶m�?      �?        ffffff�?333333�?9��8���?�q�q�?�������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�Y�Y�?;�;��?vb'vb'�?              �?�a�a�?�<��<��?F]t�E�?/�袋.�?�q�q�?9��8���?      �?                      �?              �?333333�?�������?�������?�������?      �?              �?      �?      �?                      �?�������?333333�?      �?                      �?�؉�؉�?;�;��?Cy�5��?y�5���?Nozӛ��?d!Y�B�?      �?              �?      �?�������?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?�?      �?                      �?G�<��?P���?�?p�14���?��,�?��f���?Ȥx�L�w?      �?        �{a��?�{a���? �����?8�8��?n۶m۶�?�$I�$I�?]t�E�?F]t�E�?      �?                      �?      �?              �?              �?              �?      �?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?      �?      �?        I�$I�$�?۶m۶m�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        7a~W���?�g *��?      �?        �:�r�?��دq�?к����?*�Y7�"�?              �?�������?�������?�{a���?������?              �?�������?�������?      �?        �q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        j䮟-�?e�F�t�?;ڼOq��?q�����?�c�1Ƹ?�s�9��?�ꡮ?^�^��?ffffff�?333333�?              �?      �?     ��?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?�������?�������?      �?                      �?      �?        UUUUUU�?�������?              �?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?              �?(������?6��P^C�?۶m۶m�?%I�$I��?              �?�������?ZZZZZZ�?�?�������?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?      �?      �?�m۶m��?�$I�$I�?�������?�������?      �?                      �?      �?      �?      �?                      �?              �?%I�$I��?n۶m۶�?      �?        d!Y�B�?�7��Mo�?t�E]t�?��.���?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?��8��8�?      �?      �?              �?      �?      �?              �?      �?                      �?      �?        l(�����?(������?�������?�������?              �?I�$I�$�?۶m۶m�?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�>D5hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@?         �                    �?4�5����?�           ��@                                 @E@�%W�AX�?           �z@                                   �?.��<�?)            �P@                      
             �?*;L]n�?             >@        ������������������������       �                     @                      
             �?��}*_��?             ;@                                  �Q@@�0�!��?             1@                                 �X@��S�ۿ?
             .@        	       
                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @                                   �?�z�G��?             $@                                  _@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                   @H@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                  �c@������?            �B@       ������������������������       �                     9@                                  0d@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @               /                   `@��0u���?�            �v@               *       
             �?��Q��?%             N@                                 �Z@X�EQ]N�?            �E@                                  �^@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                %                    �?�}�+r��?             C@        !       "                   �`@r�q��?             @        ������������������������       �                     @        #       $                   `j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        &       '                    �?      �?             @@       ������������������������       �                     ;@        (       )                    a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        +       ,                    �?�IєX�?             1@        ������������������������       �                      @        -       .                   `_@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        0       Y                    �?�46<�?�            �r@        1       L       	          ����?��j���?5            �T@       2       G                    �?�c�����?$            �J@       3       8                     D@ \� ���?             �H@        4       5                   g@����X�?             @        ������������������������       �                     �?        6       7                   �a@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        9       :                    �?r�q��?             E@        ������������������������       �                     $@        ;       @                    @H@     ��?             @@       <       ?                    �?�}�+r��?             3@        =       >                   0q@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        A       F                   �c@��
ц��?	             *@       B       C                   �a@      �?              @       ������������������������       �                     @        D       E                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        H       K                   0`@      �?             @        I       J                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        M       X       	          ���@*;L]n�?             >@       N       O                    �D@      �?             :@        ������������������������       �                     @        P       Q                   �a@�ՙ/�?             5@        ������������������������       �                     @        R       S                    �?և���X�?	             ,@        ������������������������       �                     @        T       W                   �r@���!pc�?             &@       U       V                   Pe@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        Z       �                   hq@�uX��?�             k@       [       j                    �?4��{���?r            @f@        \       e                    @L@Pq�����?4            @U@       ]       ^                   `l@p�|�i�?.             S@       ������������������������       �                    �D@        _       d       	             @�#-���?            �A@       `       c       
             �?�IєX�?             A@        a       b                   �\@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     =@        ������������������������       �                     �?        f       i       
             �?�����H�?             "@        g       h                    �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        k       |       
             �?��3E��?>            @W@        l       o                   ph@4���C�?            �@@        m       n                   `^@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        p       q       
             �?$��m��?             :@        ������������������������       �                      @        r       s                    �?      �?             8@        ������������������������       �                     "@        t       y                   �c@���Q��?	             .@       u       v                   0b@X�<ݚ�?             "@        ������������������������       �                      @        w       x                    `P@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        z       {                    @E@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        }       �                    �?P���Q�?'             N@        ~                           �?      �?             0@        ������������������������       �                     @        �       �                    @J@z�G�z�?             $@       ������������������������       �                     @        �       �       	          ����?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?`���i��?             F@       ������������������������       �                     C@        �       �                    a@r�q��?             @       �       �                   �_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �d@�	j*D�?            �C@       �       �                   �c@����>�?            �B@       �       �                   �`@\X��t�?             7@        ������������������������       �                     @        �       �                    @j���� �?             1@       �       �       
             �?�q�q�?	             (@        ������������������������       �                     @        �       �                    @L@�<ݚ�?             "@       ������������������������       �                     @        �       �                   @a@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        ������������������������       �                      @        �       �       
             �?l~�~��?�            0s@       �       �                   `f@�r����?�            �o@       �       �       
             �?�Zp���?�            �n@        �       �                   �a@     ��?             @@       ������������������������       �                     3@        �       �                   �b@�θ�?             *@       �       �       	             @      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @G@��Hw��?�            �j@        �       �                    �?�q�q�?             ;@       �       �                   �n@ �o_��?             9@       �       �       	          ����?     ��?             0@       �       �                   �j@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �       	              @����X�?             @        ������������������������       �                     @        �       �       	             @�q�q�?             @        ������������������������       �                     �?        �       �                    \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �       �                    �? rpa�?z            @g@        �       �       	          033�?r�q��?	             (@       �       �                    �?�C��2(�?             &@       �       �                    @I@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    c@`��F:u�?q            �e@       �       �                   P`@`k�����?n             e@        �       �                   �i@4և����?%             L@        ������������������������       �                     5@        �       �                   �^@؇���X�?            �A@        �       �                    �?�IєX�?             1@       ������������������������       �        	             ,@        �       �                    _@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    ]@�<ݚ�?             2@        �       �                    �?      �?              @       �       �                    �M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        I             \@        �       �       	             �?      �?             @        ������������������������       �                     �?        �       �                   �a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   u@      �?             $@       �       �                    g@      �?              @       �       �       	          ����?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �R@��
ц��?             J@       �       �                    k@z�J��?            �G@        �       �                    �?���y4F�?             3@       �       �                   �Y@$�q-�?	             *@       ������������������������       �                      @        �       �                   pd@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �]@      �?             @        ������������������������       �                      @        �       �                    @K@      �?             @        ������������������������       �                      @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   xr@����X�?             <@       �       �                   �\@"pc�
�?             6@        ������������������������       �                      @        �       �                   pq@ףp=
�?             4@       �       �                    �?�IєX�?	             1@       �       �                    �K@@4և���?             ,@       ������������������������       �                     &@        �       �                    �P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    d@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�   Np	�?���Gw{�?4�����?��Y>��?o�Wc"=�?IT�n��?�������?""""""�?      �?        B{	�%��?_B{	�%�?�������?ZZZZZZ�?�?�������?      �?      �?              �?      �?                      �?      �?        ffffff�?333333�?�������?UUUUUU�?              �?      �?              �?      �?      �?                      �?к����?��g�`��?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?""""""�?ffffff�?�������?qG�wĽ?w�qG�?333333�?�������?      �?                      �?(�����?�5��P�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?�������?�������?      �?                      �?�?�?      �?        �q�q�?�q�q�?      �?                      �?H�z�G�?�z�G��?�e�@	o�?o4u~�!�?�V�9�&�?:�&oe�?
^N��)�?և���X�?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?                      �?�������?UUUUUU�?      �?              �?      �?�5��P�?(�����?�������?UUUUUU�?      �?                      �?      �?        �;�;�?�؉�؉�?      �?      �?      �?              �?      �?              �?      �?                      �?      �?      �?      �?      �?              �?      �?              �?        �������?""""""�?      �?      �?              �?�<��<��?�a�a�?      �?        ۶m۶m�?�$I�$I�?      �?        t�E]t�?F]t�E�?�q�q�?�q�q�?              �?      �?              �?                      �?وlD6"�?��M�&w�?��0�9�?��x�3�?~~~~~~�?�?�k(����?^Cy�5�?      �?        �A�A�?_�_�?�?�?333333�?�������?              �?      �?              �?                      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?        '�h��&�?f�]v�e�?m��&�l�?'�l��&�?�$I�$I�?�m۶m��?      �?                      �?�N��N��?vb'vb'�?      �?              �?      �?      �?        �������?333333�?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?                      �?UUUUUU�?�������?      �?                      �?ffffff�?�������?      �?      �?      �?        �������?�������?      �?        333333�?�������?      �?                      �?F]t�E�?F]t�E�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        vb'vb'�?;�;��?�u�)�Y�?���L�?!Y�B�?��Moz��?      �?        ZZZZZZ�?�������?�������?�������?              �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?                      �?�-s�.�?�4;cS��?�?�������?�-�RM�?Az�U6�?      �?      �?              �?ى�؉��?�؉�؉�?      �?      �?      �?                      �?      �?        0x,�ն?��pB%�?UUUUUU�?UUUUUU�?�Q����?
ףp=
�?      �?      �?�q�q�?9��8���?              �?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?        �n�ᆫ?Hy�G�?UUUUUU�?�������?F]t�E�?]t�E�?�$I�$I�?۶m۶m�?      �?                      �?              �?      �?        Ȥx�L��?�u�7[��?��y��y�?�0�0�?�m۶m۶?I�$I�$�?              �?�$I�$I�?۶m۶m�?�?�?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?9��8���?      �?      �?�������?�������?              �?      �?              �?                      �?              �?      �?      �?              �?333333�?�������?      �?                      �?      �?      �?      �?      �?333333�?�������?      �?                      �?              �?      �?        �؉�؉�?�;�;�?AL� &W�?}g���Q�?(������?6��P^C�?;�;��?�؉�؉�?              �?�������?�������?              �?      �?              �?      �?      �?              �?      �?              �?      �?      �?              �?      �?        �m۶m��?�$I�$I�?/�袋.�?F]t�E�?              �?�������?�������?�?�?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���&hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK녔h��B�:         6                   Pc@({E�B��?�           ��@               #                    �?D>�Q�?`            �c@              "                   @e@�e/
�?A             [@                                  �?$	4�}�?@            �Z@                                   �O@ s�n_Y�?             J@                                 �]@X�EQ]N�?            �E@        ������������������������       �                     (@                      
             �?�חF�P�?             ?@       	                          `X@`2U0*��?             9@        
                          �S@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@                                   `@�q�q�?             @                                 @^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   a@�q�q�?             "@                                 �a@      �?              @                                 pb@���Q��?             @        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                   �M@ �Jj�G�?"            �K@       ������������������������       �                     @@                                  p`@�nkK�?             7@       ������������������������       �                     1@                !                   a@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        $       +       
             �?�q�q�?             H@       %       &                    �?      �?             @@       ������������������������       �                     7@        '       *                    �?X�<ݚ�?             "@       (       )       
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ,       5                    �P@      �?
             0@       -       .                   `Y@����X�?             ,@        ������������������������       �                      @        /       4                   �d@r�q��?             (@       0       1       	          ����?�C��2(�?             &@       ������������������������       �                      @        2       3                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        7       �                    �?N%�ξ��?p           �@        8       m       	          ����?"�ն�+�?�            `q@        9       l                     Q@�q�q��?>             X@       :       [                    �L@����X�?;            �V@       ;       J                    @G@��f/w�?(            �N@        <       G                    �?��H�}�?             9@       =       D                   �]@����X�?             5@       >       ?                    @C@�q�q�?             (@        ������������������������       �                     �?        @       C                    ]@���|���?             &@       A       B                   Hq@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        E       F       
             �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        H       I                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        K       T                    �?�����H�?             B@       L       O       
             �?�LQ�1	�?             7@        M       N                    �J@      �?             @        ������������������������       �                      @        ������������������������       �                      @        P       Q                   �c@�}�+r��?             3@       ������������������������       �        
             ,@        R       S                   @]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        U       Z                    �?$�q-�?             *@       V       Y                    @K@�����H�?             "@        W       X                    `@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        \       g                   `a@*;L]n�?             >@       ]       d                   pi@���!pc�?             6@        ^       c       
             �?X�<ݚ�?             "@       _       b                    �M@����X�?             @        `       a                    ^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        e       f                   �Y@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        h       i                    �?      �?              @        ������������������������       �                     @        j       k                    �N@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        n       �       	          ����?L�[2[
�?t            �f@        o       v                    �H@d,���O�?"            �I@        p       u                   �o@$�q-�?             *@        q       r                    �?r�q��?             @        ������������������������       �                     @        s       t                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        w       ~                   �[@�����?             C@        x       y                    �?���!pc�?             &@        ������������������������       �                     @        z       {                   l@      �?             @        ������������������������       �                      @        |       }       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @               �                   �c@PN��T'�?             ;@       �       �                    r@P���Q�?             4@       ������������������������       �        
             .@        �       �                    �L@z�G�z�?             @       ������������������������       �                     @        �       �                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     P@և���X�?             @       �       �                   �d@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �e@�Ώ��?R            ``@       �       �                   �l@P�2E��?Q            @`@        �       �                    �?��E�B��?!            �G@        �       �                   @l@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   @i@��-�=��?            �C@        �       �                   �h@�θ�?	             *@       �       �       	             �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                     L@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   0j@ ��WV�?             :@        �       �                    ]@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     .@        ������������������������       �        0            �T@        ������������������������       �                     �?        �       �                    @K@      �?�            �r@       �       �       	             @C���?t            `g@       �       �                    �?��?}�?s             g@       �       �       
             �?��Ͻ��?h            @e@        �       �                    �?և���X�?             5@       �       �                    �?p�ݯ��?             3@        ������������������������       �                      @        �       �                   �`@���|���?	             &@        ������������������������       �                     �?        �       �                    �?�z�G��?             $@        ������������������������       �                      @        �       �                   Pm@      �?              @        ������������������������       �                     @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        V            �b@        �       �                   `m@z�G�z�?             .@       �       �                   �b@�8��8��?             (@        �       �                   �i@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          pff�?�Q����?J            @\@       �       �       
             �?P��E��?0             R@        �       �                    �?^������?            �A@       �       �                   �r@�q�����?             9@       �       �                    @\X��t�?             7@       �       �                    �?������?
             .@        �       �                   @`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �_@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   Pp@      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        �       �                     P@�MI8d�?            �B@       �       �                   �a@      �?             8@        ������������������������       �                     @        �       �                     L@ҳ�wY;�?             1@        ������������������������       �                     @        �       �                   pd@�eP*L��?             &@       �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             *@        �       �                   �o@��P���?            �D@       �       �                    �?և���X�?             5@        ������������������������       �                     @        �       �                    �N@�t����?             1@       �       �       
             �?�C��2(�?             &@       ������������������������       �                     "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @l@�q�q�?             @       �       �                   �j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     4@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B�  Ac�Zb�?`yΨ�N�?vb'vb'�?b'vb'v�?	�%��о?_B{	�%�?�@�Ե�?��bEi�?;�;��?�;�;�?qG�wĽ?w�qG�?              �?��RJ)��?�Zk����?{�G�z�?���Q��?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ��)A��?k߰�k�?              �?d!Y�B�?�Mozӛ�?              �?UUUUUU�?�������?      �?                      �?      �?        �������?�������?      �?      �?              �?�q�q�?r�q��?UUUUUU�?�������?      �?                      �?      �?              �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?���)�?���ʻ��?ZMB��?S��u@7�?�������?�������?�m۶m��?�$I�$I�?XG��).�?��!XG�?{�G�z�?
ףp=
�?�m۶m��?�$I�$I�?�������?�������?              �?]t�E]�?F]t�E�?9��8���?�q�q�?      �?                      �?              �?�q�q�?�q�q�?              �?      �?              �?      �?      �?                      �?�q�q�?�q�q�?��Moz��?Y�B��?      �?      �?      �?                      �?�5��P�?(�����?      �?        �������?�������?              �?      �?        �؉�؉�?;�;��?�q�q�?�q�q�?      �?      �?              �?      �?              �?              �?        """"""�?�������?F]t�E�?t�E]t�?�q�q�?r�q��?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?        �؉�؉�?;�;��?              �?      �?              �?      �?              �?�������?�������?              �?      �?                      �?�!�!�?��{��{�?PPPPPP�?�������?;�;��?�؉�؉�?UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?^Cy�5�?Q^Cy��?F]t�E�?t�E]t�?      �?              �?      �?      �?              �?      �?      �?                      �?h/�����?&���^B�?�������?ffffff�?              �?�������?�������?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?333333�?�������?      �?                      �?              �?#����[�?^�WqBJ�?z�z��?_�^��?AL� &W�?�l�w6��?      �?      �?              �?      �?        �A�A�?}˷|˷�?�؉�؉�?ى�؉��?�q�q�?�q�q�?      �?                      �?      �?      �?              �?      �?        ;�;��?O��N���?F]t�E�?]t�E�?      �?                      �?              �?              �?      �?              �?      �?�=�����?*�Ap*�?��ׄ���?�	A����?NNNNNN�?�?�$I�$I�?۶m۶m�?^Cy�5�?Cy�5��?      �?        F]t�E�?]t�E]�?      �?        333333�?ffffff�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�8�1�s�?�c�:F�?�q�q�?r�q��?_�_��?uPuP�?���Q��?�p=
ף�?��Moz��?!Y�B�?�?wwwwww�?333333�?�������?              �?      �?        �������?�������?      �?                      �?      �?      �?      �?                      �?      �?                      �?��L���?L�Ϻ��?      �?      �?      �?        �������?�������?      �?        ]t�E�?t�E]t�?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        �����?������?۶m۶m�?�$I�$I�?      �?        �������?�������?F]t�E�?]t�E�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�EhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@=         �                    �?�r,��?�           ��@              a       	          ����?�K8c�?            z@                                 @E@&�Op��?�            �k@                      
             �?      �?'             P@       ������������������������       �                     D@                      	             �?r�q��?             8@              
                     E@�LQ�1	�?             7@               	                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                      	          ����?�X�<ݺ?
             2@                                  e@ףp=
�?             $@                                  �K@z�G�z�?             @        ������������������������       �                     @                                  �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?               R       	          pff�? �q(���?g            �c@              +                    _@��Zy�?M            @]@                                  @W@�q�q�?             B@        ������������������������       �                     @               (       	             �?      �?             @@                                  �F@�������?             >@        ������������������������       �                     �?                                   �?V�a�� �?             =@        ������������������������       �                     �?               '                   `q@�>4և��?             <@              "                   �h@PN��T'�?             ;@                !       
             �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        #       $                   l@P���Q�?
             4@       ������������������������       �                     $@        %       &       
             �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        )       *                     L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ,       A                   `q@�q�q�?8            @T@       -       :                    �L@��6}��?(            �N@       .       1       
             �?,���i�?            �D@        /       0                    �I@      �?             @        ������������������������       �                      @        ������������������������       �                      @        2       3                   �c@�L���?            �B@       ������������������������       �                     9@        4       5                   �c@      �?             (@        ������������������������       �                      @        6       9                    m@ףp=
�?             $@        7       8                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ;       >       	          ����?�G�z��?             4@       <       =                   Pd@r�q��?
             (@       ������������������������       �                     $@        ������������������������       �                      @        ?       @                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        B       Q                   xu@�G�z��?             4@       C       P       	          ����?     ��?             0@       D       I                    s@������?             .@        E       H                    s@      �?              @       F       G                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        J       K       
             �?և���X�?             @        ������������������������       �                     @        L       O                   `c@      �?             @       M       N                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        S       `                   �`@0,Tg��?             E@       T       U                    �?r�q��?             8@        ������������������������       �                     "@        V       _                    a@�r����?             .@       W       ^                    �?      �?              @       X       Y                   l@����X�?             @        ������������������������       �                     �?        Z       ]                   @_@r�q��?             @        [       \                    @I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        b       q                    �?��A� �?t             h@        c       n       
             �?*
;&���?             G@       d       g       	          ����?�˹�m��?             C@        e       f                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        h       m                   �c@�X�<ݺ?             B@        i       j       
             �?r�q��?             (@        ������������������������       �                     �?        k       l                    �?"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     8@        o       p                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        r       {       	          033�?@9G��?X            `b@        s       t                    @L@0�)AU��?%            �L@       ������������������������       �                     ?@        u       v                    _@ ��WV�?             :@       ������������������������       �                     5@        w       z                     M@z�G�z�?             @        x       y                    Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        |       �                    s@�X�<ݺ?3            �V@       }       �                    �?���(-�?+            @R@       ~       �                   @b@     �?$             P@              �       
             �?�]0��<�?"            �N@       �       �                    _@ �Jj�G�?            �K@        �       �       	          `ff@$�q-�?             *@       ������������������������       �                      @        �       �                   �p@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     E@        �       �                    �N@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �P@�t����?             1@       ������������������������       �                     .@        ������������������������       �                      @        �       �                    `@�.j�[��?�            �s@        �       �                    �?k�q��?6            @U@       �       �                    �L@Nd^����?'            �N@       �       �       
             �?�'�`d�?            �@@        �       �                    �?�q�q�?             "@       �       �                    @K@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @c@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        �       �                   p@X�Cc�?             <@       �       �       
             �?      �?             ,@       �       �                    �?�q�q�?
             (@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    a@d}h���?             ,@        �       �                   @[@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   p`@      �?             8@        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             0@        �       �       
             �?�Nx�1�?�             m@        �       �                    �?      �?/             R@        �       �                    c@�8��8��?             8@       �       �       	          ����?�nkK�?             7@       ������������������������       �                     .@        �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?�q���?              H@        ������������������������       �                     @        �       �       	          833�?�K��&�?            �E@        �       �                   0a@�8��8��?             (@        �       �                    �?z�G�z�?             @       �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?`՟�G��?             ?@       �       �                    �?�f7�z�?             =@       �       �                   @i@�G��l��?             5@        ������������������������       �                     @        �       �                   �l@j���� �?             1@        �       �       	            �?      �?              @        �       �                    `P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ]@�q�q�?	             "@        ������������������������       �                     �?        �       �       	            �?      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @       �       �                    c@      �?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ��� @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���`uӽ?h             d@       �       �                    @F��}��?\            @b@       �       �                     L@h�����?Y            �a@       ������������������������       �        N            �^@        �       �       	          ��� @�t����?             1@       �       �                   �a@      �?
             0@        ������������������������       �                      @        �       �                   ps@؇���X�?	             ,@       �       �                    �L@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    l@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �`@�r����?             .@       �       �                    �L@�8��8��?	             (@       ������������������������       �                     "@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �292ȯ�?�f����?�N��N��?O��N���?��b�#?�?��4n`�?      �?      �?              �?UUUUUU�?�������?Y�B��?��Moz��?�������?333333�?              �?      �?        �q�q�?��8��8�?�������?�������?�������?�������?              �?      �?      �?              �?      �?                      �?              �?      �?        ���c��?%w�΀�?� � �?\��[���?UUUUUU�?UUUUUU�?      �?              �?      �?�������?�������?      �?        a���{�?��{a�?      �?        �m۶m��?�$I�$I�?h/�����?&���^B�?۶m۶m�?�$I�$I�?              �?      �?        �������?ffffff�?              �?�������?�������?              �?      �?              �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?�!XG��?;ڼOq��?�����?8��18�?      �?      �?              �?      �?        }���g�?L�Ϻ��?      �?              �?      �?              �?�������?�������?      �?      �?              �?      �?              �?        �������?�������?UUUUUU�?�������?              �?      �?              �?      �?      �?                      �?�������?�������?      �?      �?�?wwwwww�?      �?      �?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?        1�0��?�y��y��?UUUUUU�?UUUUUU�?      �?        �?�������?      �?      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?              �?�LF�W>�?b6�5��?8��Moz�?���,d!�?^Cy�5�?��P^Cy�?      �?      �?      �?                      �?�q�q�?��8��8�?UUUUUU�?�������?              �?F]t�E�?/�袋.�?      �?                      �?              �?      �?      �?      �?                      �?9/���?������?p�}��?��Gp�?              �?;�;��?O��N���?              �?�������?�������?      �?      �?              �?      �?                      �?�q�q�?��8��8�?�P�B�
�?��իW��?      �?     ��?;ڼOqɠ?\2�h��?��)A��?k߰�k�?;�;��?�؉�؉�?              �?�������?�������?      �?                      �?              �?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�?<<<<<<�?              �?      �?        ��k#֥�?g@(�S��?]]]]]]�?QQQQQQ�?�u�y���?���:�?6�d�M6�?'�l��&�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?�������?UUUUUU�?              �?      �?        �m۶m��?%I�$I��?      �?      �?�������?�������?      �?              �?      �?      �?                      �?      �?        ۶m۶m�?I�$I�$�?      �?      �?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?              �?�X����?����S�?      �?      �?UUUUUU�?UUUUUU�?�Mozӛ�?d!Y�B�?      �?              �?      �?              �?      �?                      �?�������?�������?      �?        ���)k��?��)kʚ�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?              �?              �?�1�c��?�s�9��?O#,�4��?a���{�?��y��y�?1�0��?              �?�������?ZZZZZZ�?      �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?      �?      �?                      �?              �?              �?      �?      �?      �?                      �?              �?��.�?��6ͯ?��Ǐ?�?����?�m۶m��?�$I�$I�?      �?        �������?�������?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?                      �?      �?      �?              �?      �?        �������?�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ4�phG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKυ�h��B�3         v                    �?z��K���?�           ��@              M       
             �?��$����?           |@                      	          ����?���k&�?k            �g@               	                    �F@�y��*�?              M@                                   �?���Q��?             $@        ������������������������       �                     @                                  `a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        
              
             �?      �?             H@        ������������������������       �                      @                                  �X@��<b�ƥ?             G@                                   �?�C��2(�?             &@        ������������������������       �                     @                                  �W@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �A@               6                    a@B��仱�?K            �`@                     	          ����? �.�6��?-             W@                                  �p@ ��WV�?             :@       ������������������������       �                     3@                                   �L@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @               1       	          ����?����e��?            �P@              .                   @c@��6���?             E@                                 �T@     ��?             @@        ������������������������       �                     @               #                    ]@����"�?             =@               "                    �M@      �?              @                !                    �K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        $       +                   b@�G��l��?
             5@       %       &                    �E@�	j*D�?             *@        ������������������������       �                      @        '       (                    �?"pc�
�?             &@       ������������������������       �                     @        )       *                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ,       -       	          033�?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        /       0       
             �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        2       3                     O@      �?             8@       ������������������������       �        	             .@        4       5                    �O@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        7       8                   �\@��P���?            �D@        ������������������������       �                     $@        9       :                    �I@¦	^_�?             ?@        ������������������������       �                     @        ;       H                    �?��H�}�?             9@       <       G                    �?��
ц��?             *@       =       B       	          ����?���Q��?	             $@        >       ?                   `c@      �?             @        ������������������������       �                      @        @       A                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        C       D                    �?r�q��?             @        ������������������������       �                     @        E       F                   �c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        I       L                    f@r�q��?             (@       J       K       	            �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        N       g                    �?�����?�             p@        O       X                    P@b����o�?,            �R@        P       W                    �?8�Z$���?             *@       Q       R                    \@���Q��?             @        ������������������������       �                     �?        S       T                   �X@      �?             @        ������������������������       �                      @        U       V                    �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        Y       Z                   pc@��a�n`�?%             O@       ������������������������       �                    �D@        [       `                    �?����X�?             5@        \       ]                    �?      �?             @        ������������������������       �                      @        ^       _                    �E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        a       b                    @I@z�G�z�?
             .@       ������������������������       �                     $@        c       f       	          ����?���Q��?             @        d       e                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        h       u       	          ���@0�,��?q            �f@       i       t                     R@X;��?n            @f@       j       o                    d@`���i��?m             f@       k       n                   �_@����X�?H             \@        l       m                   `_@ �q�q�?             8@       ������������������������       �                     7@        ������������������������       �                     �?        ������������������������       �        8             V@        p       q                    @M@     �?%             P@       ������������������������       �        #             N@        r       s                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        w       �                    @G@�Rc���?�            �q@        x       y                   `a@p�ݯ��?             C@        ������������������������       �                     2@        z       }                   �n@�z�G��?             4@       {       |                   `e@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ~       �       	          ����?r�q��?             @               �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����?�            �n@        �       �       
             �?^������?            �A@       �       �                   @_@V�a�� �?             =@        �       �                   �`@X�Cc�?             ,@        �       �                   @_@      �?              @        ������������������������       �                     �?        �       �       	             �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?��au���?�            �j@       �       �                    @��GEI_�?v            �f@       �       �       
             �?��E�"�?u            �f@        ������������������������       �                     6@        �       �                    @K@�p=
�c�?e             d@        ������������������������       �                     I@        �       �                    �P@ףp=
�?F            �[@       �       �                   `f@,sI�v�?:            �V@       �       �                   �[@�+I�9��?9            @V@        �       �                    �O@���y4F�?             C@       �       �                    �?�t����?             A@       �       �                    �?�J�4�?             9@       �       �                    b@z�G�z�?             4@       �       �                   ph@���Q��?             $@        ������������������������       �                     @        �       �                    �M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                   �b@`'�J�?%            �I@       �       �                   �`@@�E�x�?#            �H@       ������������������������       �                     D@        �       �                   pb@�����H�?             "@       ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                   `c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?        �       �                   �X@8^s]e�?             =@        ������������������������       �                      @        �       �                    �?������?             ;@       �       �                    �?�q�q�?             5@       �       �                    �?�z�G��?             4@       �       �                    �?8�Z$���?             *@        �       �       	          ����?r�q��?             @       �       �                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �N@؇���X�?             @       �       �                    _@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @`@և���X�?             @        ������������������������       �                      @        �       �                   �]@���Q��?             @        ������������������������       �                     �?        �       �                   b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  K�ۚ��?�)|�� �?�J��*�?l�kz��?@0$[Ds�?��m�]��?GX�i��?�4�rO#�?�������?333333�?              �?�������?�������?      �?                      �?      �?      �?      �?        d!Y�B�?��7��M�?F]t�E�?]t�E�?              �?UUUUUU�?�������?              �?      �?                      �?���7G��?d\��?����7��?�B����?O��N���?;�;��?      �?        ۶m۶m�?�$I�$I�?              �?      �?        6�d�M6�?e�M6�d�?b�a��?=��<���?      �?      �?      �?        �i��F�?	�=����?      �?      �?      �?      �?              �?      �?                      �?��y��y�?1�0��?vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?      �?              �?      �?      �?                      �?      �?      �?              �?      �?        �������?�������?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�����?������?              �?�RJ)���?��Zk���?              �?
ףp=
�?{�G�z�?�;�;�?�؉�؉�?�������?333333�?      �?      �?      �?              �?      �?              �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?�������?F]t�E�?]t�E�?      �?                      �?      �?        "o���?�!oȻ?�X�%��?�6�i�?;�;��?;�;��?�������?333333�?      �?              �?      �?              �?      �?      �?              �?      �?                      �?�s�9��?�c�1Ƹ?      �?        �m۶m��?�$I�$I�?      �?      �?              �?      �?      �?              �?      �?        �������?�������?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�ݮ��?�/�Ʈ?�u�{���?�E(B�?F]t�E�?F]t�E�?n۶m۶�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?             ��?      �?      �?              �?      �?      �?                      �?              �?              �?�Q)z��?��u�	��?Cy�5��?^Cy�5�?              �?ffffff�?333333�?n۶m۶�?�$I�$I�?      �?                      �?UUUUUU�?�������?      �?      �?      �?                      �?              �?��2��?��M����?_�_��?uPuP�?a���{�?��{a�?�m۶m��?%I�$I��?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?�?�������?              �?      �?              �?        ~�	�[�?0��>���?;ڼOqɰ?�d����?����?���?              �?�������?�������?              �?�������?�������?��I��I�?l�l��?�as�ü?�3��g�?(������?6��P^C�?�?<<<<<<�?{�G�z�?�z�G��?�������?�������?�������?333333�?              �?�������?�������?      �?                      �?              �?              �?              �?      �?        �?�������?9/���?և���X�?              �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?      �?                      �?      �?        	�=����?|a���?      �?        {	�%���?B{	�%��?UUUUUU�?UUUUUU�?333333�?ffffff�?;�;��?;�;��?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?              �?      �?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJLxhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@/         n                    �?�Z���?�           ��@              9                    �K@
��x�?           �z@                                  P@T<�K<B�?�            pq@                      	          �����8����?             7@        ������������������������       �                      @                                  �_@���N8�?             5@       ������������������������       �                     "@                      
             �?�q�q�?             (@       	       
                    �?؇���X�?             @        ������������������������       �                      @                                    J@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �I@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?               .       
             �?    ���?�             p@                                  ``@�\����?+            �P@                                    F@�t����?
             1@                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@                                  �b@ڡR����?!            �H@                                    C@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@                                   �?��+��?            �B@                      	          @33�?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?                +                   �p@��>4և�?             <@       !       *                   ``@X�<ݚ�?             2@       "       %                   `]@�n_Y�K�?
             *@        #       $                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        &       )                   �d@؇���X�?             @        '       (       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ,       -                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        /       0                    �? r���?u            �g@        ������������������������       �        )             O@        1       8                   �]@      �?L             `@        2       3                   �[@�㙢�c�?             7@       ������������������������       �                     0@        4       7                   �p@և���X�?             @       5       6                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        @            @Z@        :       W       
             �?      �?`             c@       ;       >       
             �?��C"�b�?7            �T@        <       =                   @`@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        ?       P                    �?z�G�z�?/            �Q@       @       G                    �?P����?             C@        A       B                    ]@�q�q�?             "@        ������������������������       �                     @        C       F                    `P@���Q��?             @       D       E       	          `ff�?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        H       O       	          ����?>���Rp�?             =@       I       J                   @^@     ��?             0@        ������������������������       �                     @        K       L                   k@�	j*D�?	             *@        ������������������������       �                     @        M       N                   �n@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        Q       R                    �?      �?             @@       ������������������������       �                     .@        S       T                    �?�IєX�?
             1@       ������������������������       �                     (@        U       V       	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        X       ]                   @E@d}h���?)            �Q@        Y       Z                    �N@؇���X�?             @        ������������������������       �                     @        [       \                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ^       _                   @Y@؇���X�?%            �O@        ������������������������       �                     @        `       m       	             @ףp=
�?$             N@       a       b                   �a@ 	��p�?#             M@        ������������������������       �                     7@        c       h                    �?(N:!���?            �A@        d       e                   �a@�z�G��?	             $@        ������������������������       �                     �?        f       g                    s@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        i       j                   ht@`2U0*��?             9@       ������������������������       �                     4@        k       l                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        o       �                   `f@�/oD�?�            �r@       p       �                    �?h�[F���?�            `r@        q       �       
             �?     ��?             @@       r       u                    @G@>���Rp�?             =@        s       t                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        v       �                   �s@      �?             8@       w       x                   �j@�����?             5@        ������������������������       �                     @        y       z                   �k@      �?
             0@        ������������������������       �                     �?        {       �                   @`@��S�ۿ?	             .@        |                          �`@z�G�z�?             @       }       ~       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �       	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?�1����?�            `p@       �       �                    \@�kb97�?�            �l@        �       �                    �?`�Q��?             9@        ������������������������       �                     @        �       �                    �?�KM�]�?             3@       �       �                   `_@      �?	             0@       ������������������������       �                      @        �       �                    �K@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �]@�q�q�?             @        ������������������������       �                     �?        �       �                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   0c@p� V�?�            �i@       �       �                   P`@�M����?�            @i@        �       �                   �s@hA� �?0            �Q@       �       �                    \@0�,���?-            �P@        �       �                    �?$�q-�?             :@       �       �                   �^@ףp=
�?             4@        ������������������������       �                     (@        �       �                    �J@      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �X@r�q��?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �D@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        P            �`@        �       �                   �o@      �?             @        ������������������������       �                      @        �       �                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @e@�4�����?             ?@       �       �       	             �?      �?             <@        �       �                   ``@�z�G��?             $@        �       �                    @L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     @        �       �                    �?�q�q�?             "@       �       �                   �b@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �H���x�?����C�?ɲ�F�?n����s�?\�f���?��d>�;�?8��Moz�?d!Y�B�?      �?        ��y��y�?�a�a�?              �?�������?�������?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?        �������?�������?      �?                      �?      �?     ��?>����?���>��?�?<<<<<<�?      �?      �?      �?                      �?              �?����S��?����X�?UUUUUU�?UUUUUU�?              �?      �?        *�Y7�"�?�S�n�?�q�q�?�q�q�?              �?      �?        ۶m۶m�?I�$I�$�?�q�q�?r�q��?;�;��?ى�؉��?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?�������?      �?                      �?9�{n�S�?�X�0Ҏ�?      �?              �?      �?�7��Mo�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?      �?              �?      �?dp>�c�?���|��?�������?�������?      �?                      �?�������?�������?Q^Cy��?�P^Cy�?UUUUUU�?UUUUUU�?      �?        �������?333333�?      �?      �?              �?      �?              �?        GX�i���?�i��F�?      �?      �?      �?        ;�;��?vb'vb'�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?�?�?              �?�������?�������?              �?      �?        I�$I�$�?۶m۶m�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?              �?�������?�������?������?�{a���?      �?        |�W|�W�?�A�A�?ffffff�?333333�?              �?9��8���?�q�q�?      �?                      �?���Q��?{�G�z�?      �?        �������?�������?      �?                      �?              �?�옥��?�ę֞��?���+ݻ?!͎Z��?      �?      �?GX�i���?�i��F�?�������?�������?      �?                      �?      �?      �?�a�a�?=��<���?              �?      �?      �?      �?        �?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ����?J�eDP�?�cj`?�Y�	qV�?{�G�z�?��(\���?      �?        (�����?�k(���?      �?      �?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?��,�?����`�?�F�tj�?䮟-V��?_�_�?���?g��1��?Ez�rv�?;�;��?�؉�؉�?�������?�������?              �?      �?      �?      �?      �?              �?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?      �?              �?      �?        ��RJ)��?���Zk��?      �?      �?ffffff�?333333�?      �?      �?              �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?�������?333333�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW��8hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKǅ�h��B�1         N       	          ����?�r,��?�           ��@              %       
             �?����l�?�            @w@                                   �?*T7��?L            @_@                     	          833�?���tT��?7            �U@                                 �m@ ����?*            @P@       ������������������������       �                    �H@                                   �?      �?             0@               	                   �`@      �?             @        ������������������������       �                      @        
                          �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@                                   b@�G��l��?             5@                                 �g@�q�q�?
             .@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @                                   @a@�q�q�?            �C@                                  �?�G�z��?             4@                                  @C@     ��?
             0@        ������������������������       �                      @                                   �?d}h���?	             ,@        ������������������������       �                     @                                   �?�z�G��?             $@                                  �?      �?              @       ������������������������       �                     @                                   ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        !       $                    �?�KM�]�?             3@        "       #                   Pp@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        &       -                    P@4�O)��?�            �n@        '       *                    @I@և���X�?	             ,@       (       )                   `[@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        +       ,                   �Y@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        .       G                   Pb@�8h
Q��?�             m@       /       @                    �O@��<D�m�?{            �h@       0       1                   �b@`h���?v            �g@        ������������������������       �        4            @T@        2       7                    �?h�WH��?B             [@        3       6                   �c@���|���?             6@        4       5       	          @33�?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             (@        8       ?                    �? qP��B�?3            �U@        9       :                    @F@r�q��?             (@        ������������������������       �                     @        ;       >                   @d@����X�?             @       <       =                    @J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        +            �R@        A       B                    �?����X�?             @        ������������������������       �                     �?        C       D                   pa@r�q��?             @        ������������������������       �                     @        E       F                   Pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        H       I                   �b@���"͏�?            �B@        ������������������������       �                     @        J       K                   d@6YE�t�?            �@@       ������������������������       �                     .@        L       M                    �?�E��ӭ�?
             2@        ������������������������       �                     @        ������������������������       �                     *@        O       �                    �?~_d+�^�?�            �v@       P       c                    �?hu��W�?�             o@        Q       Z                    `@��Q���?             D@        R       Y                   @^@��S���?	             .@       S       T                   @]@�<ݚ�?             "@        ������������������������       �                     �?        U       X       	             �?      �?              @        V       W                   Hq@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        [       `                   �v@H%u��?             9@       \       _                   pd@���7�?             6@        ]       ^                     L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             2@        a       b                    @O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        d       �                   �c@4S)$&�?�             j@       e       p                    @G@�v�\�?~            �i@        f       o                    �?�q�q�?             8@       g       n       
             �?�㙢�c�?             7@       h       i                   �_@��s����?             5@        ������������������������       �                     (@        j       m                    b@X�<ݚ�?             "@       k       l       	             @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        q       t                   �Q@P���Q�?q            �f@        r       s                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        u       �                    �? p�/��?o            @f@        v       }       
             �?��� ��?             ?@       w       |                    X@ ��WV�?             :@        x       {                    `@؇���X�?             @        y       z       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        ~                           �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �[@P����?X            `b@        �       �                    �?�q�q�?             @       �       �                   Pl@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    _@��V9��?S            �a@        �       �                   �[@$�q-�?             *@        ������������������������       �                     @        �       �                   �\@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          033�?     ��?K             `@       ������������������������       �        (            �P@        �       �                    c@��v$���?#            �N@       ������������������������       �                      L@        �       �                   Pc@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�z1�9��?D            @\@        �       �                   �c@д>��C�?             =@       �       �       	          ����?$�q-�?             :@        �       �                   `X@؇���X�?             ,@        ������������������������       �                     �?        �       �                    �?$�q-�?             *@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �        	             (@        ������������������������       �                     @        �       �                    `@�D����?1             U@        �       �       	             �? �Cc}�?             <@        ������������������������       �                     �?        �       �                    �?�>����?             ;@        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �? �q�q�?             8@        �       �       	          `ff�?      �?              @        �       �                   �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     0@        �       �       	          ���@h�����?!             L@       �       �                   �`@0,Tg��?             E@       �       �       
             �?ܷ��?��?             =@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �K@$�q-�?             :@        ������������������������       �                     �?        �       �                   �q@`2U0*��?             9@       ������������������������       �                     2@        �       �                   �r@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�n_Y�K�?
             *@       �       �       	             �?      �?             $@       �       �                    �?r�q��?             @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�Bp  �292ȯ�?�f����?�DM4��?^v�e�]�?�~j�t��?B`��"��?�}A_�?����/��? �����? �����?              �?      �?      �?      �?      �?              �?      �?      �?      �?                      �?              �?��y��y�?1�0��?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?I�$I�$�?۶m۶m�?      �?        ffffff�?333333�?      �?      �?      �?              �?      �?              �?      �?                      �?              �?(�����?�k(���?UUUUUU�?UUUUUU�?      �?                      �?              �?���/>�?��Q���?۶m۶m�?�$I�$I�?�$I�$I�?۶m۶m�?      �?                      �?�m۶m��?�$I�$I�?              �?      �?        R��L��?m�����?��S�r
�?և���X�?�䣓�N�?p����?      �?        ��^B{	�?B{	�%��?]t�E]�?F]t�E�?�������?�������?              �?      �?              �?        ��}A�?�}A_З?�������?UUUUUU�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?      �?                      �?v�)�Y7�?*�Y7�"�?              �?'�l��&�?e�M6�d�?      �?        �q�q�?r�q��?              �?      �?        �o��.��?��T4O�?q��н?ݱ�a�E�?�������?333333�?�?�������?�q�q�?9��8���?      �?              �?      �?      �?      �?              �?      �?                      �?      �?        ���Q��?)\���(�?F]t�E�?�.�袋�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?P���?�?��	x>�?�������?�������?�������?UUUUUU�?d!Y�B�?�7��Mo�?�a�a�?z��y���?              �?�q�q�?r�q��?UUUUUU�?�������?              �?      �?              �?                      �?      �?        �������?ffffff�?      �?      �?      �?                      �?p�\��?�G?�я�?�B!��?�{����?;�;��?O��N���?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?              �?333333�?�������?      �?                      �?���+ݛ?�_��!�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?t�n���?�D�)͋�?;�;��?�؉�؉�?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?     ��?              �?;ڼOqɐ?.�u�y�?              �?�������?�������?      �?                      �?�������?�������?      �?                      �?��M�l�?6h�e�&�?a���{�?|a���?�؉�؉�?;�;��?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?      �?      �?              �?      �?              �?              �?                      �?z��y���?�0�0�?۶m۶m�?%I�$I��?      �?        h/�����?�Kh/��?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?n۶m۶�?%I�$I��?�y��y��?1�0��?��=���?a���{�?UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?;�;��?              �?���Q��?{�G�z�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ى�؉��?;�;��?      �?      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��UhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK녔h��B�:         �                    �?��}���?�           ��@                                 �`@�/<�"�?           @{@                                   @O@\�CX�?+            �Q@                                  �?lGts��?!            �K@               
                    �?�q�q�?             2@                                 �_@ףp=
�?             $@       ������������������������       �                     @               	                    `@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     @                                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �B@                                   �?      �?
             0@                                   �P@ףp=
�?             $@        ������������������������       �                     @                                   �Q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                      	             @r�q��?             @       ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               G                    �?d����?�            �v@               @       	          ����?A�b��?I            �\@              5       	          833�?v�X��?:             V@                      
             �?�0u��A�?(             N@        ������������������������       �        	             ,@        !       *                   `\@�3Ea�$�?             G@        "       #                   �b@b�2�tk�?
             2@        ������������������������       �                      @        $       )                   �[@�z�G��?             $@       %       &                   �g@���Q��?             @        ������������������������       �                     �?        '       (       	          ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        +       .                    �?@4և���?             <@        ,       -                    b@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        /       4                   pj@���N8�?             5@        0       1                    b@      �?             @        ������������������������       �                      @        2       3                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        6       7                   f@ �Cc}�?             <@        ������������������������       �                     �?        8       9                    �?�>����?             ;@        ������������������������       �                     &@        :       ;                   �[@      �?             0@        ������������������������       �                     �?        <       =       	          ����?��S�ۿ?             .@       ������������������������       �                     &@        >       ?                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        A       D                   `c@���B���?             :@       B       C                    `Q@�C��2(�?             6@       ������������������������       �                     4@        ������������������������       �                      @        E       F                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        H       o                   �`@��Pak��?�            `o@       I       V                   0k@`1�=7q�?e            �c@        J       Q                    �?��pBI�?)            @R@        K       L       	          ����?�C��2(�?             &@        ������������������������       �                      @        M       N                    �?�q�q�?             @        ������������������������       �                     �?        O       P                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        R       S       	          ����?0�z��?�?$             O@       ������������������������       �        "             N@        T       U                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        W       n       	          ��� @H��?"�?<             U@       X       e                    @L@�Zl�i��?9            @T@       Y       \                   �l@�IєX�?0             Q@        Z       [       
             �?؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        ]       d       
             �? 7���B�?)             K@        ^       c                    @�<ݚ�?             "@       _       b       	          ����?      �?              @        `       a                    @J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        !            �F@        f       m                   �p@�	j*D�?	             *@       g       h                   �Y@      �?              @        ������������������������       �                      @        i       j                    _@�q�q�?             @        ������������������������       �                     �?        k       l                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        p       �       
             �?��k=.��?E            �W@        q       x                    �?      �?             :@        r       s                    �?ףp=
�?             $@        ������������������������       �                     @        t       u                   @c@z�G�z�?             @        ������������������������       �                     @        v       w                   0l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        y       �                    �?      �?             0@       z       �                   �c@r�q��?             (@       {       |                    @z�G�z�?             $@        ������������������������       �                     @        }       ~                     N@���Q��?             @        ������������������������       �                     �?               �                   �l@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   `_@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �       	          033@����p�?4             Q@       �       �                   �c@�L#���?3            �P@        ������������������������       �                     >@        �       �                    �?������?            �B@       �       �                   xt@�t����?             A@       �       �                   �`@      �?             @@        �       �                   Pi@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �K@(;L]n�?             >@       ������������������������       �                     6@        �       �                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?��� ��?�            �r@       �       �                   �b@��Н�z�?�            p@       �       �                    �?�e)���?�            �m@        �       �                    �?�'�`d�?            �@@       �       �                   �^@���}<S�?             7@        �       �                   �[@���Q��?             @        ������������������������       �                     �?        �       �                    Z@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             2@        �       �       
             �?      �?             $@        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                     L@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   `f@�IєX�?            �i@       �       �                   @Y@ ��A�4�?}             i@        ������������������������       �                     �?        �       �                   �[@�X�� �?|             i@        �       �                    �?R���Q�?             4@       �       �                    �K@�θ�?	             *@       ������������������������       �                     @        �       �                   �p@      �?             @       �       �       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          `ff @(;L]n�?p            �f@       �       �                   �b@�nkK�?V            @a@       �       �                    �L@P�c0"�?@            @Z@       �       �                    @K@@9G��?!            �H@       ������������������������       �                    �A@        �       �                   �\@؇���X�?             ,@        �       �                   �Z@���Q��?             @       �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     L@        �       �                   �_@<���D�?            �@@       �       �       
             �? ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                    �?և���X�?             @       �       �                   `c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     E@        �       �                    @N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�z�G��?             4@        ������������������������       �                     @        �       �                   `c@      �?	             0@       �       �                    �D@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    k@��]�T��?            �D@        �       �                   pd@�����H�?             2@       �       �                    �?�IєX�?             1@       ������������������������       �                     *@        �       �                    @K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          pff�?\X��t�?             7@       �       �                   @`@r�q��?
             (@        �       �                   �^@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?���!pc�?             &@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  q��H��?��>���?��p=�?^8�߅�?��V��?=�]���?�־a�?�<%�S��?UUUUUU�?UUUUUU�?�������?�������?              �?�������?�������?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?              �?      �?      �?�������?�������?      �?              �?      �?              �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        ���}a)�?���	zZ�?�,�����?-����b�?�.�袋�?颋.���?�������?�������?              �?����7��?��,d!�?�8��8��?9��8���?      �?        333333�?ffffff�?333333�?�������?              �?      �?      �?      �?                      �?              �?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?                      �?��y��y�?�a�a�?      �?      �?      �?              �?      �?              �?      �?              �?        %I�$I��?۶m۶m�?              �?�Kh/��?h/�����?      �?              �?      �?              �?�������?�?      �?              �?      �?              �?      �?        ى�؉��?��؉���?F]t�E�?]t�E�?              �?      �?              �?      �?              �?      �?        g��1=�?��0p��?b��x�Y�?�\�:�2�?���Ǐ�?����?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        |���{�?�B!��?      �?              �?      �?              �?      �?        �<��<��?1�0��?�"e����?�����H�?�?�?۶m۶m�?�$I�$I�?              �?      �?        	�%����?h/�����?9��8���?�q�q�?      �?      �?      �?      �?              �?      �?              �?                      �?      �?        vb'vb'�?;�;��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?                      �?g���Q��?br1���?      �?      �?�������?�������?      �?        �������?�������?      �?              �?      �?              �?      �?              �?      �?UUUUUU�?�������?�������?�������?              �?�������?333333�?      �?              �?      �?      �?                      �?              �?      �?      �?              �?      �?        �������?�����Ҳ?��@���?g��1��?      �?        ��g�`��?к����?<<<<<<�?�?      �?      �?      �?      �?      �?                      �?�������?�?      �?              �?      �?              �?      �?                      �?      �?                      �?7`��c.�?��Ug��?���?����?�Ӭ����?�e��Ao�?'�l��&�?6�d�M6�?d!Y�B�?ӛ���7�?�������?333333�?              �?      �?      �?              �?      �?                      �?      �?      �?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?              �?      �?                      �?�?�?�C��x�?��`ph�?      �?        
ףp=
�?���(\��?333333�?333333�?�؉�؉�?ى�؉��?              �?      �?      �?      �?      �?              �?      �?                      �?              �?�?�������?d!Y�B�?�Mozӛ�?8�8��??�c?�c�?9/���?������?              �?�$I�$I�?۶m۶m�?�������?333333�?      �?      �?              �?      �?              �?                      �?              �?|���?|���?;�;��?O��N���?      �?                      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?333333�?ffffff�?      �?              �?      �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?jW�v%j�?KԮD�J�?�q�q�?�q�q�?�?�?              �?      �?      �?              �?      �?              �?        !Y�B�?��Moz��?�������?UUUUUU�?333333�?�������?      �?                      �?      �?        t�E]t�?F]t�E�?              �?      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��DphG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@A         �                    �?���-�g�?�           ��@              '                    �?�p�?	           0z@                                  ``@�G\�c�?(            @P@              	                     D@���Q��?            �A@                      	          `ff�?r�q��?             @                                  �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        
                           �?8^s]e�?             =@                                  �?R���Q�?             4@                                 �s@�t����?             1@       ������������������������       �        
             .@        ������������������������       �                      @                                   ^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                      	             �?�q�q�?             "@                      	          @33�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               "       
             �?z�G�z�?             >@              !                    �?HP�s��?             9@                                  �o@r�q��?             (@                                  �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �M@ףp=
�?             $@        ������������������������       �                     @                       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             *@        #       &                    �?z�G�z�?             @       $       %                   d@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        (       M                    �G@�:�B��?�             v@        )       B       	             �?�q�q�?)            @Q@       *       /                   �k@      �?             D@        +       .                   �[@      �?	             0@        ,       -                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        0       7                    @F@�q�q�?             8@        1       6                    ]@և���X�?             @       2       5                    @E@���Q��?             @       3       4                   Hq@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        8       ;                    �?�t����?             1@        9       :       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        <       A                   @`@$�q-�?             *@        =       >                   �\@؇���X�?             @        ������������������������       �                      @        ?       @       
             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        C       D                   �Z@ܷ��?��?             =@        ������������������������       �                     �?        E       L       	             �?@4և���?             <@        F       G                    @F@؇���X�?             ,@       ������������������������       �                     @        H       K       
             �?����X�?             @       I       J                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             ,@        N       q       	          033�?|�����?�            �q@        O       ^                    �J@���!pc�?:             V@        P       [                   pc@      �?             8@       Q       R                   �X@     ��?             0@        ������������������������       �                     @        S       Z       	          ����?8�Z$���?
             *@       T       U                   �_@z�G�z�?             $@        ������������������������       �                     �?        V       W                   �a@�����H�?             "@       ������������������������       �                     @        X       Y       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        \       ]                   �`@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        _       l       	          833�?     ��?*             P@       `       k                   �d@ףp=
�?              I@       a       d                   �Y@Hm_!'1�?            �H@        b       c       
             �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        e       f       
             �?�7��?            �C@       ������������������������       �                     <@        g       j       	          ����?"pc�
�?	             &@       h       i                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        m       p                    �?      �?
             ,@       n       o                    V@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        r       �                    c@�����?~            �h@       s       �                   �_@8��"s�?u            �f@        t       {                    �?r�q��?             B@       u       v                   0`@$�q-�?             :@       ������������������������       �                     4@        w       z                    �?�q�q�?             @       x       y                    a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        |       �                    �?���Q��?             $@       }       ~                   `U@      �?              @        ������������������������       �                      @               �                    p@�q�q�?             @        ������������������������       �                      @        �       �                   �p@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �R@P����?]            `b@       �       �                    c@@��t��?[             b@       �       �                    Y@`�LVXz�?@            �X@        �       �                    �M@�X�<ݺ?             2@        �       �                   0a@      �?              @        �       �                    �K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        5            @T@        �       �                   �l@�nkK�?             G@        �       �                     M@ףp=
�?             4@       ������������������������       �                     ,@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?d}h���?	             ,@        �       �                     P@      �?             @       �       �       	          ���@      �?             @       �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?�b��-8�?�            �s@        �       �                    �?     ��?U             `@       �       �                    �?��}E��?8            �T@        �       �                   hq@؇���X�?             <@       �       �                    �?�8��8��?             8@        �       �                   �k@      �?              @        ������������������������       �                     @        �       �                     L@�q�q�?             @        ������������������������       �                     �?        �       �                   p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �g@      �?
             0@        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �       	          `ff�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   e@���|���?'            �K@       �       �                    @�7����?#            �G@       �       �       	          ����?���"͏�?            �B@        �       �                    �?��S�ۿ?             .@        �       �                   �\@r�q��?             @        ������������������������       �                     @        �       �                   @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �c@���|���?             6@       �       �                   �`@�z�G��?             4@       �       �       
             �?���Q��?             .@        �       �       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?
             (@        �       �                     D@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �F@�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �b@���Q��?             $@        ������������������������       �                     @        �       �                   �c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �L@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @Y@:	��ʵ�?            �F@        ������������������������       �                      @        �       �                   �e@(L���?            �E@       �       �                   �`@��-�=��?            �C@       �       �       
             �?(;L]n�?             >@        ������������������������       �                     @        �       �                   p`@ ��WV�?             :@        �       �                   @_@@4և���?             ,@       ������������������������       �                     "@        �       �       	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             (@        �       �                   �l@�q�q�?             "@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    @F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �M@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �                          �Q@���ͫt�?s            `g@       �             	          `ff�?hl �&�?r             g@       �       �                    �?�ګ���?n            `f@        ������������������������       �        .            �R@        �                           �?P�c0"�?@            @Z@       �       �                    @L@p�C��?8            �V@       ������������������������       �        +            @Q@        �       �                    �?�C��2(�?             6@       �       �                   @a@8�Z$���?	             *@        ������������������������       �                     @        �       �                   0b@�q�q�?             @        ������������������������       �                     �?        �       �                   ps@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     ,@                                `U@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��hb�BP  lk�w��?J��	.�?��^Wۓ�?S(*	[�?[��Z���?S+�R+��?333333�?�������?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?|a���?	�=����?333333�?333333�?<<<<<<�?�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�������?�������?{�G�z�?q=
ףp�?UUUUUU�?�������?      �?      �?              �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?      �?      �?                      �?      �?        �pR���?�c+����?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?      �?      �?                      �?              �?UUUUUU�?�������?�$I�$I�?۶m۶m�?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        <<<<<<�?�?      �?      �?              �?      �?        �؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?              �?        a���{�?��=���?      �?        �$I�$I�?n۶m۶�?�$I�$I�?۶m۶m�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�	�Z��?��Q)z��?t�E]t�?F]t�E�?      �?      �?      �?      �?              �?;�;��?;�;��?�������?�������?              �?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?              �?      �?�������?�������?9/���?Y�Cc�?�������?�������?              �?      �?        �A�A�?��[��[�?              �?F]t�E�?/�袋.�?      �?      �?              �?      �?                      �?      �?              �?      �?ffffff�?333333�?              �?      �?                      �?�����?/,FBi��?�k�g��?E���Y@�?UUUUUU�?�������?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?�������?333333�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?���+ݛ?�_��!�?��RA�/�?*h���V�?[�R�֯�?�~�@��?�q�q�?��8��8�?      �?      �?      �?      �?              �?      �?                      �?              �?              �?d!Y�B�?�Mozӛ�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?        ۶m۶m�?I�$I�$�?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?�u]�u]�?QEQE�?      �?      �?�7�:���?��ˊ��?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        F]t�E�?]t�E]�?G}g����?]AL� &�?*�Y7�"�?v�)�Y7�?�?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?F]t�E�?]t�E]�?333333�?ffffff�?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?                      �?      �?        �������?333333�?              �?�������?�������?      �?                      �?      �?      �?      �?                      �?l�l��?��O��O�?      �?        w�qG��?⎸#��?�A�A�?}˷|˷�?�?�������?              �?;�;��?O��N���?�$I�$I�?n۶m۶�?              �?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?                      �?              �?      �?      �?              �?      �?        v^��u�?��/G��?ozӛ���?Y�B��?!�R"x��?�7Ck��?      �?        ?�c?�c�?8�8��?��K��K�?h�h��?      �?        ]t�E�?F]t�E�?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?              �?        �������?�������?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ%�[6hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hK
hyK�hzh)h,K ��h.��R�(KK���h��B�/         L                   p`@P��]��?�           ��@               !       	          pff�?���m/��?�            �t@                                  �a@��~�a�?P             `@                                   �?д>��C�?$             M@                                  �?�:�^���?            �F@                                  �?PN��T'�?             ;@                                 �[@������?	             1@                                   �?և���X�?             @       	       
                   �Z@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                  �_@ףp=
�?             $@       ������������������������       �                     @                      
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     2@                                   [@��
ц��?             *@       ������������������������       �                     @        ������������������������       �                     @                                   �?R_u^|�?,            �Q@                     
             �?�2�o�U�?!            �K@                                    F@�X�<ݺ?	             2@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                    �B@                                   xp@      �?             0@                     	          ����?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        "       K                   �z@b �57�?�            �i@       #       4       	          ����?(���h�?            �i@        $       -                    �L@b�h�d.�?            �A@        %       &                    �?�q�q�?             .@        ������������������������       �                     @        '       (                   �_@r�q��?	             (@       ������������������������       �                      @        )       ,                    b@      �?             @       *       +                   �n@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        .       3                    @M@P���Q�?             4@        /       2                    �?؇���X�?             @        0       1                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        5       <                    \@h�|�6�?i            @e@        6       7                    �?z�G�z�?             .@        ������������������������       �                      @        8       ;                    �?$�q-�?
             *@        9       :                   `_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        =       J                   Xp@ ���l��?^            `c@       >       G                   P`@ ��WV�?@             Z@       ?       D                   0p@` A�c̭?>             Y@       @       C                   �e@��K2��?<            �W@        A       B                   Pe@�?�|�?            �B@       ������������������������       �                     B@        ������������������������       �                     �?        ������������������������       �        #            �L@        E       F                   �^@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        H       I                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �I@        ������������������������       �                     �?        M       �                    �?��d��?           �x@        N       k       
             �?�lg����?m            �e@       O       Z                    �?B�1V���?>            @X@        P       Q                   �^@���!pc�?            �@@        ������������������������       �                     @        R       S                    a@д>��C�?             =@        ������������������������       �                     (@        T       U                   `a@�t����?             1@        ������������������������       �                     @        V       Y       	          ����?؇���X�?	             ,@        W       X                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        [       j                    �?     ��?)             P@       \       ]                   �`@8�Z$���?            �C@        ������������������������       �                     �?        ^       i                    �M@�?�'�@�?             C@       _       d                    q@���B���?             :@       `       a                   �m@��S�ۿ?             .@        ������������������������       �                      @        b       c                   @n@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        e       f                   �b@���|���?             &@        ������������������������       �                     @        g       h                    @D@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     9@        l       y       	          833�?.�W����?/            �R@       m       r                    �?     ��?             H@        n       q                    p@�q�q�?             (@       o       p                   `h@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        s       t                    �?�X�<ݺ?             B@       ������������������������       �                     =@        u       v                   �c@����X�?             @        ������������������������       �                     @        w       x                   �d@      �?             @       ������������������������       �                      @        ������������������������       �                      @        z                            P@��}*_��?             ;@       {       ~                    �?��+7��?             7@       |       }                   0l@���Q��?             .@        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �K@�y!>�K�?�            `l@       �       �       
             �?������?j             d@        �       �                   Ph@�q�q�?            �F@        �       �                    �?����X�?             ,@       �       �                    �?"pc�
�?             &@        ������������������������       �                     �?        �       �                   �b@ףp=
�?             $@        �       �                    K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?�חF�P�?             ?@        �       �                   �m@���Q��?             $@        �       �                   �`@r�q��?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @���N8�?             5@       ������������������������       �                     1@        �       �                    a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        M             ]@        �       �       	          ����?�eP*L��?*            �P@       �       �                    �M@��Zy�?            �C@        �       �       
             �?b�2�tk�?             2@        ������������������������       �                     �?        �       �                    �?ҳ�wY;�?             1@       �       �                    @      �?             0@       �       �                    �L@      �?	             (@       �       �                   �q@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �O@����X�?             5@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `j@�n_Y�K�?             *@        ������������������������       �                     @        �       �                   �c@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                     P@l��
I��?             ;@       �       �                    �N@     ��?             0@       �       �                    b@"pc�
�?	             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �h6n���?���� ��?����'t�?R�����?4�9c��?�9cΘ�?|a���?a���{�?l�l��?}�'}�'�?h/�����?&���^B�?�?xxxxxx�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?      �?      �?              �?      �?                      �?              �?�؉�؉�?�;�;�?              �?      �?        �@�6�?2~�ԓ��?־a��?�S�<%��?�q�q�?��8��8�?      �?                      �?      �?              �?      �?      �?      �?              �?      �?                      �?�H%�e�?��VC��?<��;�?��߁��?_�_��?;��:���?UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?ffffff�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?�?�������?�������?�������?      �?        ;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?mЦm�?-��,�?;�;��?O��N���?���Q��?
ףp=
�?W�+�Ʌ?��Q�٨�?к����?*�Y7�"�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?                      �?      �?        �3�τ?�?�=`���?�}A_��?}A_��?��4l7��?���$2�?t�E]t�?F]t�E�?      �?        |a���?a���{�?              �?�������?�������?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?      �?;�;��?;�;��?      �?        y�5���?������?ى�؉��?��؉���?�?�������?              �?�$I�$I�?۶m۶m�?      �?                      �?F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?贁N��?0��b�/�?      �?      �?�������?�������?�m۶m��?�$I�$I�?              �?      �?                      �?��8��8�?�q�q�?      �?        �m۶m��?�$I�$I�?      �?              �?      �?              �?      �?        B{	�%��?_B{	�%�?Y�B��?zӛ����?�������?333333�?              �?      �?                      �?      �?        *�����?Y[�;���?c��*��?�싨�ٷ?UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?F]t�E�?/�袋.�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �Zk����?��RJ)��?333333�?�������?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?      �?      �?              �?      �?                      �?��y��y�?�a�a�?      �?              �?      �?              �?      �?              �?        ]t�E�?t�E]t�?� � �?\��[���?9��8���?�8��8��?      �?        �������?�������?      �?      �?      �?      �?      �?      �?              �?      �?              �?                      �?              �?�m۶m��?�$I�$I�?      �?      �?              �?      �?        ;�;��?ى�؉��?              �?�������?�������?      �?                      �?h/�����?Lh/����?      �?      �?F]t�E�?/�袋.�?              �?      �?              �?        F]t�E�?]t�E�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�	3 hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKǅ�h��B�1         .                    �?�[��N�?�           ��@                      	          `ff�?�.�+��?e            �e@              
                    �?<����??            �W@               	                   Pb@�θ�?             :@                                   N@���N8�?             5@       ������������������������       �        
             1@                                   @P@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �?��.N"Ҭ?0            @Q@                                   `@�r����?             .@       ������������������������       �                     @                                  �e@�<ݚ�?             "@        ������������������������       �                     @                                   �I@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        (             K@               +                   �c@�o;����?&            �S@              *                    `P@�ɞ`s�?            �N@              #                    @K@      �?             L@                                  �?�f7�z�?             =@                                  �H@@�0�!��?	             1@       ������������������������       �                     (@                      
             �?���Q��?             @                                  `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                   �b@      �?             (@       ������������������������       �                      @        !       "                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        $       )                    @M@�>����?             ;@        %       (                    �?z�G�z�?             $@       &       '                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     @        ,       -                    �?�����H�?             2@        ������������������������       �                      @        ������������������������       �                     0@        /       �       
             �?��~V��?f           ��@       0       }                   f@������?�             v@       1       P       	          ����?�s���?�            �u@        2       9                   �_@�L"��?D            �Z@       3       4                   @l@����˵�?&            �M@       ������������������������       �                     �I@        5       6                    �?      �?              @        ������������������������       �                     @        7       8                    _@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        :       ;                    @D@�q�q�?             H@        ������������������������       �                     $@        <       =                     E@p�ݯ��?             C@        ������������������������       �                     @        >       ?                    @J@">�֕�?            �A@        ������������������������       �                     @        @       G       	          833�?��>4և�?             <@       A       B                    @��S�ۿ?	             .@       ������������������������       �                     "@        C       F                    �?r�q��?             @       D       E                     P@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        H       I                    X@�θ�?             *@        ������������������������       �                     �?        J       O                     M@r�q��?             (@        K       L                    _@���Q��?             @        ������������������������       �                      @        M       N                   Pj@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        Q       |                    �R@ 1�/Gu�?�            �m@       R       ]                    �F@��!Dϸ?�            `m@        S       V                   �Z@��<b���?             7@        T       U                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        W       X                    �?�S����?             3@        ������������������������       �                      @        Y       Z                   �_@�IєX�?             1@        ������������������������       �                     "@        [       \                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ^       c                   @Z@ ���X�?�            �j@        _       `                   `X@z�G�z�?             @        ������������������������       �                     @        a       b                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        d       i                    �?��.N"Ҭ?�            �i@       e       f                   hr@�=
ףp�?c             d@       ������������������������       �        T             a@        g       h                   �r@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        j       w                   pb@�*/�8V�?             �G@       k       l                   0b@��p\�?            �D@       ������������������������       �                     ;@        m       n       	          `ff�?d}h���?             ,@        ������������������������       �                     @        o       v                   �`@�q�q�?             "@       p       q                    �?      �?             @        ������������������������       �                      @        r       u                    \@      �?             @        s       t       	          `ff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        x       y                   c@�q�q�?             @        ������������������������       �                     �?        z       {                    �Q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ~                           @D@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?j�*�'�?�            �i@        �       �                    �?��:��?8            @V@       �       �                    �?�D��?!            �H@       �       �                    �L@^H���+�?            �B@       �       �                    �?      �?             <@        �       �                   �^@      �?              @        ������������������������       �                      @        �       �                   pe@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �I@ףp=
�?             4@       ������������������������       �        	             (@        �       �                   @`@      �?              @        ������������������������       �                     �?        �       �                   �^@؇���X�?             @       ������������������������       �                     @        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   Xs@�q�q�?             "@       �       �                   P`@      �?              @        ������������������������       �                     @        �       �                   �c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �d@�G�z�?             D@       �       �                     O@����>�?            �B@       �       �                    �H@X�Cc�?             <@        ������������������������       �                     @        �       �       	             �?�eP*L��?             6@        �       �                   �b@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �\@�	j*D�?             *@       �       �                    �?X�<ݚ�?             "@       �       �                    @N@�q�q�?             @       �       �       	             �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                    @L@��-�=��?M            @]@       �       �                    �?��4+̰�??            @X@        �       �                     H@z�G�z�?             $@       ������������������������       �                     @        �       �                   �]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   pf@���E�?9            �U@       ������������������������       �        3            �S@        �       �       	          433�?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �L@�G�z��?             4@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?�q�q�?             .@       ������������������������       �                     "@        �       �                   Pb@r�q��?             @       ������������������������       �                     @        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�Bp  B~�9�J�?�@c�Z�?�f��o�?�2)^ �?���%N�?�X�0Ҏ�?ى�؉��?�؉�؉�?��y��y�?�a�a�?      �?              �?      �?              �?      �?                      �?�3J���?ہ�v`��?�������?�?      �?        9��8���?�q�q�?      �?              �?      �?      �?                      �?      �?        ��	�Z�?�#{���?&C��6��?mާ�d�?      �?      �?a���{�?O#,�4��?�������?ZZZZZZ�?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?              �?      �?              �?      �?        h/�����?�Kh/��?�������?�������?      �?      �?      �?                      �?              �?              �?      �?        �q�q�?�q�q�?              �?      �?        B�A��?_�_��?��)����?���%Ƨ�?�qG��?G�w��?���~!V�?��L�w��?��/���?W'u_�?              �?      �?      �?              �?333333�?�������?              �?      �?        �������?�������?              �?Cy�5��?^Cy�5�?      �?        �A�A�?_�_��?              �?I�$I�$�?۶m۶m�?�?�������?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        (�X�>�?��v��?5���	%�?-�!c�]�?��Moz��?��,d!�?      �?      �?              �?      �?        ^Cy�5�?(������?      �?        �?�?              �?      �?      �?      �?                      �?�	�[��?e�Cj���?�������?�������?              �?      �?      �?              �?      �?        ہ�v`��?�3J���?������y?�������?              �?UUUUUU�?�������?      �?                      �?m�w6�;�?r1����?��+Q��?�]�ڕ��?              �?۶m۶m�?I�$I�$�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?        333333�?�������?              �?      �?        WC���?R�yY�'�?�x�3��?�as���?������??4և���?L�Ϻ��?�g�`�|�?      �?      �?      �?      �?      �?        UUUUUU�?�������?              �?      �?        �������?�������?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?���L�?�u�)�Y�?�m۶m��?%I�$I��?              �?]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?                      �?;�;��?vb'vb'�?�q�q�?r�q��?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        }˷|˷�?�A�A�?_\����? tT����?�������?�������?      �?              �?      �?              �?      �?        m��֡�?Ȥx�L��?      �?              �?      �?      �?                      �?�������?�������?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKŅ�h��B@1         v       
             �?�_y���?�           ��@              M                    �?T:�:w��?	           �x@                                  �g@�xO��(�?g             c@                                  �^@4և����?$             L@               
                    T@r�q��?             2@              	                    �?$�q-�?	             *@                                   �K@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   �F@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                   @Q@�}�+r��?             C@                                  �?��?^�k�?            �A@       ������������������������       �                     8@                                  �`@�C��2(�?             &@                                   �?�q�q�?             @                                  �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               .                    �?�d�~V��?C            @X@               -                   {@�q�q�?             E@                                 �Z@�(�Tw��?            �C@        ������������������������       �                     @                                   @i@�<ݚ�?             B@        ������������������������       �                      @        !       "       
             �?@�0�!��?             A@        ������������������������       �                     @        #       $                   �_@�n`���?             ?@        ������������������������       �                     (@        %       (                    b@�����?             3@        &       '                   0a@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        )       *                    �?8�Z$���?	             *@        ������������������������       �                     @        +       ,       	             �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        /       <                   �o@ؓ��M{�?'            �K@       0       1                    �?�z�G��?             >@        ������������������������       �                     &@        2       ;       	          ��� @�\��N��?             3@       3       4                   �\@�q�q�?             .@        ������������������������       �                     @        5       8                   �a@r�q��?
             (@        6       7                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        9       :                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        =       @                    �J@���Q��?             9@        >       ?                    d@      �?              @        ������������������������       �                     @        ������������������������       �                     @        A       F                    �?�t����?             1@        B       C                    �?      �?              @        ������������������������       �                     @        D       E                   Xr@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        G       L                   0b@�����H�?             "@        H       I                     @      �?             @        ������������������������       �                      @        J       K                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        N       Q                    Z@p�����?�             n@        O       P                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        R       o                   �b@0�����?�            �m@       S       l                   `f@0���|�?�             l@       T       e                   �s@ �й���?�            `k@       U       ^                    �?`�LVXz�?�            �h@       V       ]                    �D@�Ŗ�Pw�?\            @a@        W       \                    `@@4և���?
             ,@        X       Y       
             �?z�G�z�?             @        ������������������������       �                     �?        Z       [                   `U@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        R             _@        _       d                    �J@ �.�?Ƞ?(             N@        `       a                    �I@r�q��?             @        ������������������������       �                     @        b       c                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        $             K@        f       k                   ``@���N8�?             5@        g       h                    �?z�G�z�?             @        ������������������������       �                     �?        i       j                    @L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             0@        m       n       	          ����?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        p       q       	          433�?؇���X�?	             ,@        ������������������������       �                     �?        r       u                    �?$�q-�?             *@        s       t                    @H@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        w       �                   @E@H�V�e��?�            @u@        x       �                    �?t/*�?            �G@        y       z                   �\@���|���?             6@        ������������������������       �                      @        {       �                    �?�z�G��?
             4@        |       �                   �d@      �?             $@       }       ~                    �?����X�?             @        ������������������������       �                     @               �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @b@ףp=
�?             $@       ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@        �       �                    �?ؓFl:8�?�            Pr@        �       �                    �L@`�Q��?/            �R@       �       �       	             @z�G�z�?#            �K@       �       �                    `@8�Z$���?"             J@       �       �                     K@��a�n`�?             ?@       �       �                    �?�X����?             6@        ������������������������       �                     @        �       �                   �a@j���� �?             1@        ������������������������       �                     @        �       �                    n@���|���?
             &@       �       �       	          ����?      �?              @       �       �                    ]@և���X�?             @       �       �                   @[@���Q��?             @        ������������������������       �                     �?        �       �                   d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �e@���N8�?             5@       ������������������������       �                     3@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��Q��?             4@        �       �                   �l@      �?             (@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @N@      �?              @        ������������������������       �                     @        �       �                    _@z�G�z�?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   ``@��6�.ӯ?�            @k@       ������������������������       �        N            �^@        �       �                    �?�8��8N�?5             X@       �       �                     L@��`qM|�?,            �T@       ������������������������       �                     �O@        �       �                    c@z�G�z�?             4@        ������������������������       �                     $@        �       �                    d@���Q��?             $@        ������������������������       �                      @        �       �                    �M@      �?              @       �       �                    �L@      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�θ�?	             *@       �       �       	          hff @���!pc�?             &@       �       �                   xs@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  V�.�#��?աh6n��?>�]X���?����^�?�?�?��?6��5���?�m۶m۶?I�$I�$�?UUUUUU�?�������?;�;��?�؉�؉�?UUUUUU�?�������?              �?      �?                      �?�������?333333�?      �?                      �?(�����?�5��P�?�A�A�?_�_��?              �?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �,O"Ӱ�?�i�n�'�?UUUUUU�?UUUUUU�?� � �?�o��o��?      �?        �q�q�?9��8���?      �?        �������?ZZZZZZ�?              �?�c�1��?�9�s��?              �?^Cy�5�?Q^Cy��?UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        	� O	�?�־a��?ffffff�?333333�?      �?        y�5���?�5��P�?UUUUUU�?UUUUUU�?              �?�������?UUUUUU�?      �?      �?              �?      �?        �������?�������?      �?                      �?              �?�������?333333�?      �?      �?              �?      �?        �������?�������?      �?      �?      �?        �������?�������?              �?      �?        �q�q�?�q�q�?      �?      �?              �?      �?      �?      �?                      �?              �?$�$��?���?      �?      �?      �?                      �?M�[��?��'�W2�?߼�xV4�?*;L]n�?����?����Ǐ�?[�R�֯�?�~�@��?ہ�v`�}?��?���?�$I�$I�?n۶m۶�?�������?�������?              �?      �?      �?              �?      �?                      �?              �?�?wwwwww�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�a�a�?��y��y�?�������?�������?              �?      �?      �?              �?      �?                      �?UUUUUU�?�������?      �?                      �?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?iiiiii�?ZZZZZZ�?W�+���?�;����?F]t�E�?]t�E]�?      �?        333333�?ffffff�?      �?      �?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?                      �?�������?�������?              �?      �?      �?              �?      �?                      �?ܴE��?Y���?��(\���?{�G�z�?�������?�������?;�;��?;�;��?�c�1��?�s�9��?�E]t��?]t�E]�?      �?        �������?ZZZZZZ�?      �?        F]t�E�?]t�E]�?      �?      �?�$I�$I�?۶m۶m�?�������?333333�?      �?              �?      �?              �?      �?              �?                      �?              �?      �?        ��y��y�?�a�a�?      �?              �?      �?              �?      �?                      �?ffffff�?�������?      �?      �?      �?                      �?      �?      �?              �?�������?�������?              �?      �?      �?              �?      �?        ���A���?��p�?      �?        �������?�������?�@	o4u�?��k���?      �?        �������?�������?      �?        333333�?�������?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ى�؉��?�؉�؉�?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?                      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��~hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKɅ�h��B@2         v                    �?���w���?�           ��@              K       
             �?`�Q��?            |@                      	          ����?���|���?j             f@                      
             �?���B���?             J@        ������������������������       �                     @                                   �?      �?             H@                                   Z@X�<ݚ�?             "@        ������������������������       �                     @        	       
                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �]@�7��?            �C@        ������������������������       �                     $@                                  @^@ 	��p�?             =@                                  �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �? ��WV�?             :@                                  �E@���N8�?             5@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             2@        ������������������������       �                     @               *                    �?V{q֛w�?K             _@               )                   �a@      �?%             P@                                   ]@�g�y��?             ?@                                   �M@�8��8��?             (@                                    L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        !       (                   `s@���y4F�?             3@       "       #                   @Y@r�q��?             2@        ������������������������       �                      @        $       '                    �?      �?
             0@        %       &       
             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                    �@@        +       <                   Hp@d��0u��?&             N@       ,       -                    �G@d}h���?             E@        ������������������������       �                     &@        .       /                    �?¦	^_�?             ?@        ������������������������       �                     @        0       5       	          033�?      �?             8@        1       2                    �K@      �?              @       ������������������������       �                     @        3       4                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        6       ;                    @      �?
             0@       7       :                   `d@և���X�?             ,@       8       9                   �`@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        =       >       
             �?�E��ӭ�?             2@        ������������������������       �                     �?        ?       @       	          ����?������?
             1@        ������������������������       �                     @        A       J                    �L@���|���?             &@       B       I                    @L@�q�q�?             @       C       D                   �b@      �?             @        ������������������������       �                     �?        E       H                     G@�q�q�?             @       F       G       	              @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        L       u       	          `ff@��)��g�?�             q@       M       t                   0e@,7���v�?�            �p@       N       e                    �?���PXY�?�            `j@        O       V                    �?�q�q�?%             N@        P       U                    q@�n_Y�K�?             *@       Q       R                   �a@����X�?             @        ������������������������       �                     @        S       T       	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        W       d                   �_@�*/�8V�?            �G@       X       Y                   @E@���|���?            �@@        ������������������������       �                     @        Z       [                     I@�<ݚ�?             ;@        ������������������������       �                     $@        \       _                    �J@ҳ�wY;�?             1@        ]       ^                   �l@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        `       c       	          ����?ףp=
�?             $@       a       b                   �[@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        f       m       	          pff�?������?\            �b@       g       h                    @L@؀���˲?O            ``@       ������������������������       �        C            @[@        i       j                   �b@�GN�z�?             6@       ������������������������       �                     0@        k       l       	          ����?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        n       s                    j@z�G�z�?             4@        o       p                    d@�q�q�?             @        ������������������������       �                      @        q       r                   �h@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �        '             N@        ������������������������       �                     @        w       �                    �?�������?�            �q@        x       �                   �u@��e�B��?            �I@       y       |                    �G@F�����?            �F@        z       {                   �b@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        }       �                    �?����X�?            �A@       ~       �       
             �?д>��C�?             =@              �                   `^@$�q-�?             :@        �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �                     M@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     4@        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?�/�T�?�             m@       �       �                    �?�'݊U�?X            �`@       �       �                    @K@�HP��a�?E            @[@        �       �       
             �?@9G��?            �H@       �       �                   �_@ qP��B�?            �E@        ������������������������       �                     8@        �       �                   pb@�}�+r��?             3@       ������������������������       �                     1@        �       �                    c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?d��0u��?'             N@       �       �                     P@��i#[�?             E@       �       �       	          hff�?|��?���?             ;@        �       �       	          ����?؇���X�?             @       �       �                    �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �l@��Q��?             4@        �       �                    Y@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        
             .@        ������������������������       �                     2@        �       �       
             �?� �	��?             9@       �       �                   `i@�z�G��?             4@        �       �                   �`@ףp=
�?             $@       ������������������������       �                     @        �       �                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	             �?      �?             $@        ������������������������       �                     @        �       �                    �?����X�?             @       �       �       	             �?���Q��?             @        ������������������������       �                     �?        �       �                   m@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �Z@�FVQ&�?C            �X@        ������������������������       �                      @        �       �                   8p@��8�$>�?B            @X@       ������������������������       �        '             M@        �       �                    c@��-�=��?            �C@       �       �                     R@�X�<ݺ?             B@       �       �                   �_@��?^�k�?            �A@        �       �       
             �?z�G�z�?             @        ������������������������       �                     �?        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                     �?        �       �                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  @��"z�?౏��B�?��(\���?{�G�z�?F]t�E�?]t�E]�?ى�؉��?��؉���?      �?              �?      �?�q�q�?r�q��?              �?�������?�������?      �?                      �?�A�A�?��[��[�?              �?�{a���?������?UUUUUU�?UUUUUU�?      �?                      �?;�;��?O��N���?�a�a�?��y��y�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�{����?B!��?      �?      �?�B!��?��{���?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?6��P^C�?(������?�������?UUUUUU�?              �?      �?      �?�������?�������?              �?      �?              �?                      �?              �?DDDDDD�?wwwwww�?I�$I�$�?۶m۶m�?      �?        ��Zk���?�RJ)���?      �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?              �?r�q��?�q�q�?      �?        �?xxxxxx�?              �?F]t�E�?]t�E]�?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?/�#EC�?������?2�]��?�wo�e�?Z�����?�6����?UUUUUU�?UUUUUU�?ى�؉��?;�;��?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?              �?�٨�l��?AL� &W�?]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?        �������?�������?�$I�$I�?�m۶m��?              �?      �?        �������?�������?�������?�������?              �?      �?              �?              �?        �^x/��?�z=��?h�T��?�i��?      �?        �袋.��?]t�E�?      �?        UUUUUU�?�������?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?                      �?=�]���?�9�h���?�������?�������?؂-؂-�?�>�>��?ffffff�?333333�?              �?      �?        �$I�$I�?�m۶m��?|a���?a���{�?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?        �������?UUUUUU�?      �?                      �?      �?        ����S��?Y����?��[���?����?���[��?������?9/���?������?�}A_З?��}A�?              �?(�����?�5��P�?              �?      �?      �?      �?                      �?UUUUUU�?�������?              �?      �?        �������?�?�<��<��?�a�a�?	�%����?{	�%���?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        ffffff�?�������?ffffff�?333333�?              �?      �?                      �?              �?              �?)\���(�?�Q����?333333�?ffffff�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?�m۶m��?�$I�$I�?333333�?�������?      �?              �?      �?      �?                      �?      �?              �?        |���?>����?      �?        ����?�Q�/��?              �?�A�A�?}˷|˷�?�q�q�?��8��8�?�A�A�?_�_��?�������?�������?              �?      �?      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@0         f                    �?({E�B��?�           ��@              +       	          ����?fD1�n�?           �x@                      
             �?��t�?e            �a@                                  �g@$�Z����?2             S@       ������������������������       �                    �C@                      	          833�?V������?            �B@                                  �?�>����?             ;@        ������������������������       �        	             ,@        	       
                   �b@8�Z$���?	             *@       ������������������������       �                     &@        ������������������������       �                      @                                   b@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                                  @E@@i��M��?3            @P@                                   �?؇���X�?             @                      	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �b@�BbΊ�?-             M@                                  �?XB���?             =@                                  �j@z�G�z�?             @                                   ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     8@               "                    �?l��[B��?             =@                                  �q@�����H�?             "@       ������������������������       �                     @                !                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        #       *                   �d@��Q��?             4@       $       %                    @J@@4և���?	             ,@       ������������������������       �                     @        &       )                    �?؇���X�?             @       '       (                    �K@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ,       c                    �R@�Z�)��?�            �o@       -       R       
             �?���+[��?�            `o@       .       7                   `\@���8�?�            �k@        /       0                    �?����X�?             5@        ������������������������       �                      @        1       2                   �R@���y4F�?             3@        ������������������������       �                      @        3       6                   Pk@���|���?             &@        4       5                   @a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        8       M                   �x@8be��|�?{             i@       9       F                   Pr@ E59|�?w             h@       :       E                    �?��z*�o�?`            �c@       ;       <                    @M@�T�~~4�?E            @]@       ������������������������       �        '            @S@        =       @                    �?P���Q�?             D@        >       ?                   P`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        A       D                    �M@��?^�k�?            �A@        B       C                   �`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @@        ������������������������       �                     E@        G       H                   �r@��hJ,�?             A@        ������������������������       �                     @        I       J                   �u@(;L]n�?             >@       ������������������������       �                     4@        K       L                   �e@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        N       Q       	          ����?      �?              @       O       P                    �H@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        S       ^                    �?J�8���?             =@       T       ]                    c@�G�z��?             4@       U       V                   �e@������?             .@        ������������������������       �                      @        W       \                    �?8�Z$���?	             *@        X       Y                   0l@      �?             @        ������������������������       �                     �?        Z       [       	            �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        _       b                    �?�����H�?             "@        `       a                    @F@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        d       e                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        g       ~                    `@�0��;�?�            0u@        h       }       
             �?�s��:��?0             S@       i       p       	          `ff�?���B���?!             J@        j       o                   �^@���7�?             6@        k       n                    �?؇���X�?             @       l       m                   `X@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        q       x                    �?�z�G��?             >@        r       w                    @P@�q�q�?             "@       s       t                    �?      �?             @        ������������������������       �                      @        u       v                    Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        y       z                   �s@؇���X�?             5@       ������������������������       �                     0@        {       |                   `c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     8@               �       	          ���@Θ	���?�            pp@       �       �                    @@�g8���?�            `o@       �       �       
             �?@��xQ�?�            �l@        �       �                    �G@�2�o�U�?'            �K@        ������������������������       �                     0@        �       �                   �p@��Zy�?            �C@       �       �                    �?���>4��?             <@        �       �                   pe@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             5@        �       �                   l@�q�q�?             @        ������������������������       �                     �?        �       �       	          433�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?�E��ӭ�?             2@        ������������������������       �                     �?        �       �                   �k@������?             1@        ������������������������       �                     @        �       �                    �M@�	j*D�?             *@       �       �                   �Z@z�G�z�?             $@        ������������������������       �                     �?        �       �                   �b@�����H�?             "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          `ff�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        �       �       	            �?�ً�q��?j            �e@       �       �                    �?��V9��?X            �a@        �       �                    �?      �?             0@       �       �                   0m@ףp=
�?             $@        �       �                    �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �t@ >��@�?L            @_@       ������������������������       �        J            �^@        �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          pff�?     ��?             @@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     <@        �       �                    �?
;&����?             7@       �       �                    �?     ��?             0@        ������������������������       �                     @        �       �                   �\@�q�q�?	             (@        ������������������������       �                     @        �       �                    �N@      �?              @       �       �       
             �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     O@r�q��?	             (@       ������������������������       �                     $@        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  Ac�Zb�?`yΨ�N�?ל�b8�?�XE_�1�?d-C���?Ni^����?l(�����?�5��P^�?              �?o0E>��?�g�`�|�?h/�����?�Kh/��?              �?;�;��?;�;��?              �?      �?        �������?�������?      �?                      �?�Z��Z��?�J��J��?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?�{a��?���=��?GX�i���?�{a���?�������?�������?      �?      �?      �?                      �?      �?              �?        ���=��?GX�i���?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ffffff�?�������?�$I�$I�?n۶m۶�?              �?�$I�$I�?۶m۶m�?UUUUUU�?�������?      �?                      �?              �?      �?        O���t:�?��b�X�?�';r���?���Ɏ�?�9	ą��?��~G���?�$I�$I�?�m۶m��?      �?        (������?6��P^C�?              �?F]t�E�?]t�E]�?�������?�������?      �?                      �?              �?t��2�?)��|�?�?��葢?!�~���?��N�?|mĺ���?���??�s?�s�?              �?�������?ffffff�?�������?�������?      �?                      �?�A�A�?_�_��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?KKKKKK�?      �?        �?�������?              �?�������?�������?              �?      �?              �?      �?�������?�������?              �?      �?                      �?|a���?�rO#,��?�������?�������?�?wwwwww�?      �?        ;�;��?;�;��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �q�q�?�q�q�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �~#���?���i<�?�k(���?��k(��?ى�؉��?��؉���?F]t�E�?�.�袋�?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?              �?333333�?ffffff�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?333333�?�������?      �?                      �?      �?        )�I�y��?\�Nj�?/�*�S��?D�Tw�V�?��b:���?:��,���?־a��?�S�<%��?      �?        � � �?\��[���?n۶m۶�?I�$I�$�?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?r�q��?�q�q�?      �?        �?xxxxxx�?              �?;�;��?vb'vb'�?�������?�������?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?/�袋.�?F]t�E�?      �?                      �?�6��<�?�'�j��?�D�)͋�?t�n���?      �?      �?�������?�������?      �?      �?      �?                      �?      �?              �?        X9��v��?����Mb�?      �?              �?      �?      �?                      �?      �?      �?      �?      �?              �?      �?              �?        �Mozӛ�?Y�B��?      �?      �?      �?        �������?�������?      �?              �?      �?UUUUUU�?�������?              �?      �?              �?                      �?UUUUUU�?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�DhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKŅ�h��B@1         �       
             �?&I,|-��?�           ��@              !                    �?;6��?           �y@                                   �J@և���X�?-            �Q@                                  �t@x�����?            �C@              
                    �?�MI8d�?            �B@                                   �?     ��?             0@        ������������������������       �                      @               	                   �s@      �?              @       ������������������������       �                     @        ������������������������       �                     @                      	          ����?���N8�?             5@       ������������������������       �                     &@                      	          033�?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @                                   `@¦	^_�?             ?@                                   �?�eP*L��?             &@        ������������������������       �                     @                      	            @����X�?             @       ������������������������       �                     @        ������������������������       �                      @                                    @M@z�G�z�?             4@                                   �?���Q��?             $@                                 pd@և���X�?             @                                 @q@z�G�z�?             @        ������������������������       �                      @                                  �q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             $@        "       E                   @l@�8��_��?�            pu@       #       0                   pa@=QcG��?x            �g@       $       )       
             �?@��8��?Z             b@        %       (                    �?�C��2(�?             6@        &       '                   @\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        *       +                   `\@ ��7��?K            �^@       ������������������������       �        '             Q@        ,       -                    �Q@@3����?$             K@       ������������������������       �        "            �I@        .       /       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        1       :                    �?�������?             F@       2       9                   �b@ 	��p�?             =@        3       4                   @a@z�G�z�?             $@        ������������������������       �                     @        5       8                   h@�q�q�?             @        6       7                   Pb@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     3@        ;       B                    �?��S���?             .@       <       A                    b@�z�G��?             $@        =       @                   �a@      �?             @        >       ?                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        C       D                   j@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        F       G                   �l@xG�"��?`            `c@        ������������������������       �                     @        H       c                    �?X��S���?^             c@        I       b                   �e@�+��<��?            �E@       J       _                   �r@�q�q�?             B@       K       ^       	          ���@r֛w���?             ?@       L       W                   �b@V�a�� �?             =@       M       N                    `@�q�q�?
             .@        ������������������������       �                     @        O       P                   @_@      �?             $@        ������������������������       �                     @        Q       R                    �N@����X�?             @        ������������������������       �                      @        S       V                   �b@���Q��?             @       T       U                   Pn@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        X       Y                   �d@@4և���?	             ,@        ������������������������       �                      @        Z       ]                   �d@r�q��?             @        [       \                   `m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        `       a       	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        d       i                   �[@�~i��?C            @[@        e       h                   �m@      �?              @        f       g                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        j       �                    c@ܴD��?>            @Y@       k       x                    �?�8��8N�?;             X@       l       w                    \@����!p�?4             V@        m       r                   �[@$G$n��?            �B@       n       q                   �p@      �?             @@        o       p                   (p@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             8@        s       t                   �p@z�G�z�?             @        ������������������������       �                      @        u       v                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        "            �I@        y       z                    �L@      �?              @        ������������������������       �                      @        {       ~                    �?�q�q�?             @       |       }                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               �                   0`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���Q��?             @       �       �       	          033@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�l8ɠ��?�            t@        �       �                    @N@�a�O�?;            @X@       ������������������������       �        3            @U@        �       �                   �s@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                    c@���X�?�             l@        �       �                    �?������?             A@       �       �                    �?X�<ݚ�?             2@        ������������������������       �                     �?        �       �                   0a@��.k���?             1@        �       �                    �?�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?      �?              @       �       �                    [@���Q��?             @        ������������������������       �                     �?        �       �                    @G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             0@        �       �                    @O@�"�q��?}            �g@       �       �                    �?\-��p�?r            �e@        �       �                   �l@Z��Yo��?$             O@        �       �                   �^@��2(&�?             6@        ������������������������       �                     $@        �       �                    �I@      �?
             (@        ������������������������       �                     @        �       �                   pc@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   ``@      �?             D@       �       �                   �a@��+7��?             7@        ������������������������       �                     @        �       �                    �?�X�<ݺ?             2@        ������������������������       �                     @        �       �                    �K@�8��8��?             (@       �       �                   �[@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	          pff�?@�0�!��?
             1@       ������������������������       �        	             ,@        ������������������������       �                     @        �       �                    �L@����X�?N             \@       ������������������������       �        D            �W@        �       �       	          833@�X�<ݺ?
             2@       ������������������������       �        	             1@        ������������������������       �                     �?        �       �                     P@      �?             0@        ������������������������       �                     @        �       �                    �?�q�q�?             "@       �       �                   Pp@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �"z?+�?���B`��?B�[\��?p��(V�?�$I�$I�?۶m۶m�?��o��o�?�A�A�?��L���?L�Ϻ��?      �?      �?      �?              �?      �?              �?      �?        ��y��y�?�a�a�?      �?        �������?�������?              �?      �?                      �?�RJ)���?��Zk���?]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?      �?                      �?�������?�������?�������?333333�?�$I�$I�?۶m۶m�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?��xҊ*�?��aK]��?AL� &W�?x6�;��?UUUUUU�?UUUUUU�?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?;ڼOqɀ?��:ڼ�?              �?h/�����?���Kh�?              �?UUUUUU�?UUUUUU�?              �?      �?        /�袋.�?t�E]t�?�{a���?������?�������?�������?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�?333333�?ffffff�?      �?      �?      �?      �?              �?      �?              �?                      �?�������?�������?      �?                      �?=���?������?      �?        ������?��P^Cy�?w�qG�?w�qG��?UUUUUU�?UUUUUU�?�B!��?���{��?a���{�?��{a�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        �$I�$I�?�m۶m��?              �?�������?333333�?      �?      �?      �?                      �?      �?        �$I�$I�?n۶m۶�?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?        �������?�������?              �?      �?              �?        ��A��.�?��w� z�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?z��~�X�?�(0���?�������?�������?]t�E�?/�袋.�?���L�?к����?      �?      �?      �?      �?              �?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?              �?      �?        333333�?�������?      �?      �?      �?                      �?              �?���C��?����R�? tT����?����?      �?        UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?I�$I�$�?�?xxxxxx�?�q�q�?r�q��?              �?�?�������?�q�q�?9��8���?      �?              �?      �?      �?      �?      �?                      �?              �?      �?      �?333333�?�������?              �?      �?      �?              �?      �?              �?                      �?a�+F�?|n�S���?a����?�{a���?!�B!�?���{��?��.���?t�E]t�?      �?              �?      �?      �?              �?      �?      �?                      �?      �?      �?Y�B��?zӛ����?      �?        �q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?                      �?              �?ZZZZZZ�?�������?      �?                      �?n۶m۶�?�$I�$I�?      �?        ��8��8�?�q�q�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �t�bub�G+     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���MhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@-         p       
             �?&sCA�?�           ��@              M                    �?�ދ���?           0{@                      	          ����?T#k߂�?l             e@                      
             �?�U�:��?!            �M@        ������������������������       �                     �?                                    P@ 	��p�?              M@                                 pe@ ��WV�?             J@                                  ]@@��8��?             H@        	                          @f@�8��8��?             (@       
                           �?r�q��?             @                                   �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     B@                                  f@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �a@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               "       	             �?�ϡz�?K            �[@                      	          ����?�LQ�1	�?             7@                                  �?      �?             0@                                   �?r�q��?             @        ������������������������       �                     �?                                  �[@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                !                   �`@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        #       4                    �?JyK���?9            �U@       $       )       	          ����?�q��/��?             G@        %       &                   �V@���Q��?             @        ������������������������       �                      @        '       (                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        *       1                    `Q@������?            �D@       +       0       	          ����?P�Lt�<�?             C@        ,       /                    �?      �?             @       -       .                   `]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        2       3       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        5       B                   �`@�>$�*��?            �D@        6       A                    �?և���X�?             5@       7       8                    �?��.k���?             1@        ������������������������       �                     @        9       :                   �K@�q�q�?             (@        ������������������������       �                      @        ;       @       	          033@z�G�z�?             $@       <       ?       	          ����?�����H�?             "@        =       >                   �r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        C       D                    �?�z�G��?             4@        ������������������������       �                     @        E       F                    T@@�0�!��?             1@        ������������������������       �                     �?        G       L       	          ���@      �?
             0@       H       K                    @K@��S�ۿ?	             .@        I       J                   �d@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        N       i                   �_@���}��?�            �p@       O       f       	          ����?�qE��E�?g            �d@        P       Q                   �i@�7�QJW�?-            �R@        ������������������������       �                     B@        R       S                   �[@�q�q�?            �C@        ������������������������       �                      @        T       Y                   @_@V������?            �B@        U       V                    Z@$�q-�?             *@       ������������������������       �                     "@        W       X                    \@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       c                    s@�q�q�?             8@       [       ^                   pm@�E��ӭ�?             2@        \       ]       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        _       `                    @O@�8��8��?             (@       ������������������������       �                     "@        a       b                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        d       e                    w@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        g       h                    �R@�x�E~�?:            @V@       ������������������������       �        9            �U@        ������������������������       �                      @        j       o       	          hff�?�K}��?B            �Y@        k       n                   �a@�8��8��?             (@       l       m                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        ;            �V@        q       �                    �?�㙢�c�?�            �r@       r       {                    �?0����?�            �o@        s       t                   s@�zvܰ?4             V@       ������������������������       �        +             R@        u       z       	          ����?     ��?	             0@       v       y                    �?�z�G��?             $@        w       x                    �L@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        |       �                    �?X�;�^o�?n            �d@       }       �       	            �?�:�^���?[            �`@       ~       �                    �O@��?^�k�?I            @Z@              �                   Pb@�K}��?G            �Y@       ������������������������       �        A            �V@        �       �                    @L@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          033@�z�G��?             >@       �       �                    �M@      �?             <@        �       �                   �_@�q�q�?             (@        ������������������������       �                     @        �       �                    @L@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                      @        �       �                    �?�z�G��?             >@        �       �       	          ����?և���X�?             ,@       �       �                    �?      �?              @        ������������������������       �                     @        �       �                    @E@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �Q@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        �       �                    �?�û��|�?             G@       �       �                    @N@�\��N��?             C@       �       �       	             �?��}*_��?             ;@        �       �                    p@؇���X�?             ,@       �       �                   `c@"pc�
�?             &@        ������������������������       �                      @        �       �                   �Y@�q�q�?             @        ������������������������       �                     �?        �       �                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�n_Y�K�?	             *@        ������������������������       �                      @        �       �                    c@���!pc�?             &@       �       �                    Z@�����H�?             "@        �       �                   �X@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�C��2(�?             &@        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �ۚ��?*|�� q�?�P-
��?ث��J�?&�q-�?m��1G��?�pR�屵?�A�I�?      �?        �{a���?������?;�;��?O��N���?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        yJ���?~��7�}�?��Moz��?Y�B��?      �?      �?�������?UUUUUU�?      �?        �������?�������?              �?      �?              �?        �m۶m��?�$I�$I�?      �?                      �?p��f��?Ȥx�L��?��Mozӻ?�B����?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?������?p>�cp�?(�����?���k(�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �����?�18���?�$I�$I�?۶m۶m�?�?�������?              �?UUUUUU�?UUUUUU�?              �?�������?�������?�q�q�?�q�q�?      �?      �?              �?      �?              �?                      �?      �?        333333�?ffffff�?      �?        �������?ZZZZZZ�?      �?              �?      �?�?�������?      �?      �?              �?      �?                      �?      �?        ���̮?4�τ?�?jW�v%j�?�+Q��?0��b�/�?t�@�t�?              �?UUUUUU�?UUUUUU�?      �?        o0E>��?�g�`�|�?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?�������?�������?r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?      �?                      �?p�\��?����G�?              �?      �?        �?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?�7��Mo�?d!Y�B�?[
����?'���H�?颋.���?t�E]t�?      �?              �?      �?ffffff�?333333�?�������?333333�?      �?                      �?      �?              �?        �־a��?J��yJ�?}�'}�'�?l�l��?_�_��?�A�A�?�������?�?      �?        ]t�E�?F]t�E�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ffffff�?333333�?      �?      �?�������?�������?              �?�m۶m��?�$I�$I�?      �?                      �?      �?                      �?ffffff�?333333�?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?              �?      �?                      �?      �?      �?      �?                      �?��,d!�?8��Moz�?�5��P�?y�5���?_B{	�%�?B{	�%��?۶m۶m�?�$I�$I�?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        ى�؉��?;�;��?      �?        t�E]t�?F]t�E�?�q�q�?�q�q�?�������?�������?              �?      �?                      �?      �?        F]t�E�?]t�E�?              �?UUUUUU�?�������?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ9M�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKŅ�h��B@1         p                    �?F���?��?�           ��@                                 @E@,���8k�?           0z@                      
             �?z�G�z�?,            �R@              	                    �? �h�7W�?             �J@                                  �?�(\����?             D@                                   �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     >@        
                           �?8�Z$���?             *@        ������������������������       �                     �?                      	          `ff@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?                                   �N@�eP*L��?             6@                                  \@X�Cc�?             ,@        ������������������������       �                     @                                   �?ףp=
�?             $@                                  �`@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               C       
             �?������?�            �u@               :                   @a@��|��L�?F            �\@              7                    �?R_u^|�?.            �Q@              $       	          ����?���Q��?*            @P@                !                   pe@�8��8��?	             (@       ������������������������       �                     $@        "       #                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       6       	          ��� @�#ʆA��?!            �J@       &       '                    �?���c�H�?            �H@        ������������������������       �                     9@        (       1                    �?r�q��?             8@       )       0                   r@�q�q�?
             .@       *       /                    �I@�C��2(�?             &@        +       ,                   �m@�q�q�?             @        ������������������������       �                     �?        -       .                   8p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        2       3                   �_@�����H�?             "@       ������������������������       �                     @        4       5                    �M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        8       9                    �M@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ;       <                    �N@�������?             F@        ������������������������       �                     1@        =       B                    @�q�q�?             ;@       >       A       	          ����?؇���X�?             5@        ?       @                    �?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        D       S                    �?��Q���?�            �l@        E       H                   �k@�X����?             F@        F       G       	          ����?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        I       J                     L@     ��?             @@        ������������������������       �                     &@        K       R                   �u@�ՙ/�?
             5@       L       Q                    �?�E��ӭ�?             2@       M       N                    d@      �?             $@        ������������������������       �                     @        O       P                    r@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        T       U                   @i@@-�_ .�?x             g@        ������������������������       �        "            �I@        V       Y                   pi@t�e�í�?V            �`@        W       X                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       m                    @����?T            @`@       [       ^                   @Y@/����?P            �^@        \       ]                    c@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        _       f       	            �?���<_�?M            �]@       `       a                    �?�K}��?B            �Y@       ������������������������       �        0             S@        b       c                     O@ ��WV�?             :@       ������������������������       �                     8@        d       e                    s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        g       h                    �?      �?             0@        ������������������������       �                      @        i       l                    �M@      �?              @        j       k                    r@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        n       o                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        q       �       
             �?b�h�d.�?�            �s@       r       �                    �R@���� �?�             q@       s       �                    \@��GXT1�?�            �p@        t       y                    �?X�<ݚ�?             ;@        u       x                    �K@�<ݚ�?             "@        v       w                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        z                           �?�E��ӭ�?
             2@       {       |                    �?������?	             1@       ������������������������       �                     (@        }       ~       	             �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `f@{*�?�?�             n@       �       �                   �b@��F�M�?�            �l@       �       �                   Pe@ଡ଼R�?�             j@        ������������������������       �        '            �O@        �       �                   �e@�c!�^�?a            @b@        ������������������������       �                     �?        �       �                   xp@����=O�?`             b@       �       �       	          ����?XI�~�?7            @S@        �       �                    �?؇���X�?             <@        ������������������������       �                     $@        �       �       	          ����?�<ݚ�?             2@        ������������������������       �                     @        �       �                    @K@�q�q�?             (@        ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@@�E�x�?%            �H@       ������������������������       �        "            �F@        �       �                    b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @^@ ��ʻ��?)             Q@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        %            �O@        �       �                   Pc@����X�?             5@        �       �       	          033�?�q�q�?             @       �       �       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�r����?             .@        �       �       	          ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �^@"pc�
�?             &@        ������������������������       �                     @        �       �                   �`@����X�?             @        ������������������������       �                     �?        �       �                    @N@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�+��<��?!            �E@        ������������������������       �                     "@        �       �       	          ����?�ʻ����?             A@        �       �                    �?�E��ӭ�?             2@       �       �                     N@�	j*D�?
             *@       ������������������������       �                     "@        ������������������������       �                     @        �       �                    a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             0@       ������������������������       �        	             $@        �       �       	          033�?�q�q�?             @        ������������������������       �                      @        �       �                    ^@      �?             @        ������������������������       �                     �?        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  ,�U�)�?js���?�6"�M��?���d��?�������?�������?"5�x+��?��sHM0�?�������?333333�?�������?�������?              �?      �?                      �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        t�E]t�?]t�E�?�m۶m��?%I�$I��?      �?        �������?�������?�������?�������?              �?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?������?0�����?���9E�?&��~]�?�@�6�?2~�ԓ��?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        e�Cj���?5�x+��?4և����?/�����?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?        �q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?�������?              �?      �?        /�袋.�?t�E]t�?              �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        j�$s��?����fԺ?�E]t��?]t�E]�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?        �a�a�?�<��<��?r�q��?�q�q�?      �?      �?      �?        �$I�$I�?�m۶m��?      �?                      �?              �?      �?        S�n0E�?к����?      �?        �1����?�rv��?      �?      �?      �?                      �?n�Fn�F�?�����?��/����?�M!Ф?333333�?�������?      �?                      �?+����/�?��/���?�������?�?      �?        O��N���?;�;��?      �?              �?      �?      �?                      �?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �m۶m��?�$I�$I�?      �?                      �?_�_��?;��:���?<<<<<<�?xxxxxx�?��ʹ?���¯��?�q�q�?r�q��?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        r�q��?�q�q�?�?xxxxxx�?              �?�������?�������?      �?                      �?      �?         �ޯ?���?�(�j�?�~]R�0�?wo���%�?	��u���?              �?Ĉ#F��?t�Ν;w�?      �?        ��RA�/�?U��K��?V~B����?5�wL��?�$I�$I�?۶m۶m�?              �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        9/���?և���X�?              �?      �?      �?      �?                      �?�?�������?�������?�������?      �?                      �?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?                      �?      �?      �?              �?      �?        w�qG��?w�qG�?      �?        <<<<<<�?�������?�q�q�?r�q��?vb'vb'�?;�;��?      �?                      �?�������?�������?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJpVhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK߅�h��B�7         f       	          ����?T8���?�           ��@                                 @E@����?�            pw@                                  �[@�k�'7��?$            �L@                                   �? �q�q�?             8@              
                    �?���N8�?             5@                                 �W@$�q-�?             *@       ������������������������       �                     @               	                   �^@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                      
             �?���!pc�?            �@@       ������������������������       �                     3@                                   �?X�Cc�?             ,@                                   �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @                                    E@      �?              @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               Y                    �? {��e�?�            �s@              0                    �?\|/��j�?�            �p@               %                    �?p�eU}�??            �Y@               "                    s@ȵHPS!�?             :@              !                   �_@P���Q�?             4@                                   �K@؇���X�?             @       ������������������������       �                     @                                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        #       $                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        &       '                   �Z@`<)�+�?0            @S@        ������������������������       �                     �?        (       /                    �?P�Lt�<�?/             S@        )       .                    �?r�q��?             (@       *       -       	          ����?�<ݚ�?             "@       +       ,       
             �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        (             P@        1       H       
             �?���z��?k             d@        2       9                     J@�%^�?            �E@        3       4       	          ����?���N8�?             5@       ������������������������       �                     0@        5       8                    �H@z�G�z�?             @       6       7                   8p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        :       ;       
             �?�eP*L��?             6@        ������������������������       �                      @        <       C                    �?���Q��?             4@       =       >       	          ����?���|���?             &@        ������������������������       �                      @        ?       @                    �?�<ݚ�?             "@       ������������������������       �                     @        A       B                    _@      �?             @        ������������������������       �                      @        ������������������������       �                      @        D       G                    �?�����H�?             "@       E       F       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        I       N                   `\@ ,��-�?M            �]@        J       K                    �?�q�q�?	             .@        ������������������������       �                     @        L       M                     I@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        O       T                    @L@ f^8���?D            �Y@       P       S                    �?�E�����?;            �V@        Q       R                    �B@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        5            �S@        U       X                    _@8�Z$���?	             *@        V       W       	          @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        Z       a                    �?��}*_��?             K@       [       \       
             �?�%^�?            �E@        ������������������������       �                     $@        ]       `                    �?Pa�	�?            �@@        ^       _                   @r@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     8@        b       e                    �J@"pc�
�?             &@        c       d       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        g       �                    �?*����?�            pv@       h       {                    �?�+Ĺ+�?�             o@        i       p                    �?>a�����?             �I@        j       k                   �]@ҳ�wY;�?
             1@        ������������������������       �                     @        l       m                   �a@      �?             (@        ������������������������       �                     @        n       o                   pc@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        q       z                    �?�IєX�?             A@        r       w                    �?      �?
             0@       s       t       
             �?$�q-�?             *@       ������������������������       �                     &@        u       v                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        x       y                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        |              	          033�? ���v��?z            �h@        }       ~       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?P�2E��?x            `h@       �       �                    `R@��
���?Y            �b@       �       �                   @^@PL��V�?W            �b@        �       �       	          `ff�?$�q-�?             :@        ������������������������       �                      @        �       �                   p`@�����H�?
             2@       �       �                    �?�IєX�?	             1@       �       �       	          ����?@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    c@ ��7��?G            �^@       ������������������������       �        B            �\@        �       �                     L@؇���X�?             @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �J@�����H�?            �F@        �       �                   Pm@�θ�?             *@        ������������������������       �                     @        �       �                    @G@      �?              @        ������������������������       �                     �?        �       �                   �`@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?      �?             @@       �       �                    �M@�����H�?             2@       �       �                    �?؇���X�?	             ,@       �       �                   �Y@�<ݚ�?             "@       �       �                    @M@؇���X�?             @        ������������������������       �                     @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        �       �                   �`@�eP*L��?B            �[@        �       �                   P`@������?            �B@        �       �                    `@�	j*D�?
             *@       �       �                    @O@z�G�z�?             $@       ������������������������       �                     @        �       �       	          `ff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    [@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        �       �                    �?��T���?*            @R@        �       �                   �c@�����H�?             ;@        �       �                   0c@�θ�?             *@       �       �       
             �?�C��2(�?             &@        �       �                   @q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             ,@        �       �                    �?
;&����?             G@       �       �                   0c@����e��?            �@@       �       �                   `p@�\��N��?
             3@       �       �                    �?�	j*D�?             *@        ������������������������       �                     @        �       �                   m@X�<ݚ�?             "@       �       �                    b@�q�q�?             @        ������������������������       �                      @        �       �                    @F@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    b@d}h���?	             ,@       �       �                   0r@8�Z$���?             *@       �       �       	             �?�8��8��?             (@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          ����?�	j*D�?             *@        ������������������������       �                      @        �       �                    b@z�G�z�?             @        ������������������������       �                     @        �       �                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  6n����?�� ���?�o�2z[�? ��I�?Lg1��t�?-����b�?UUUUUU�?�������?�a�a�?��y��y�?;�;��?�؉�؉�?              �?UUUUUU�?�������?      �?                      �?              �?              �?t�E]t�?F]t�E�?              �?%I�$I��?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ~�	�[�?
�[���?m��&�l�?N6�d�M�?(�J��"�?��VCӭ?��N��N�?�؉�؉�?ffffff�?�������?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        S{����?��O���?              �?���k(�?(�����?�������?UUUUUU�?9��8���?�q�q�?�m۶m��?�$I�$I�?              �?      �?              �?              �?              �?        \|r��?��6��?�}A_�?�}A_��?�a�a�?��y��y�?              �?�������?�������?      �?      �?      �?                      �?              �?]t�E�?t�E]t�?      �?        �������?333333�?]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?�������?�������?              �?      �?                      �?[4���?'u_[�?UUUUUU�?UUUUUU�?              �?�������?UUUUUU�?      �?                      �?H%�e�?��VCӝ?P��O���?l�l��?]t�E�?F]t�E�?              �?      �?              �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?        _B{	�%�?B{	�%��?�}A_��?�}A_�?              �?|���?|���?�q�q�?�q�q�?      �?                      �?      �?        F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?����>�?Ɔ��O��?���ˊ��?(፦ί�?�?�������?�������?�������?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?        �?�?      �?      �?;�;��?�؉�؉�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?1ogH�۩?�y;Cb�?UUUUUU�?UUUUUU�?              �?      �?        z�z��?_�^��?O贁N�?&�X�%�?L�Ϻ��?�u�)�Y�?;�;��?�؉�؉�?              �?�q�q�?�q�q�?�?�?�$I�$I�?n۶m۶�?      �?                      �?              �?      �?        ;ڼOqɀ?��:ڼ�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�q�q�?�q�q�?�؉�؉�?ى�؉��?              �?      �?      �?      �?        �$I�$I�?�m۶m��?      �?                      �?      �?      �?�q�q�?�q�q�?�$I�$I�?۶m۶m�?�q�q�?9��8���?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?      �?              �?      �?                      �?              �?              �?]t�E�?t�E]t�?к����?��g�`��?;�;��?vb'vb'�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�B�
*�?�z��ի�?�q�q�?�q�q�?ى�؉��?�؉�؉�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �Mozӛ�?Y�B��?6�d�M6�?e�M6�d�?y�5���?�5��P�?;�;��?vb'vb'�?              �?�q�q�?r�q��?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?        ۶m۶m�?I�$I�$�?;�;��?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?        vb'vb'�?;�;��?      �?        �������?�������?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�,         P       	          ����?6������?�           ��@              E                    �?�^�����?�            0x@                                  �?��vn[+�?�            �s@                                    L@X;��?:            @V@       ������������������������       �        ,            �P@                                  @_@�LQ�1	�?             7@        ������������������������       �                     $@               	                   �`@�θ�?	             *@        ������������������������       �                      @        
                          �c@�C��2(�?             &@        ������������������������       �                     @                                   �?      �?             @                                  �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @               &       
             �?�+̸�?�            `l@                      	          ����?8�Z$���?*            @P@                                  �?�1�`jg�?$            �K@       ������������������������       �                    �B@                                   j@r�q��?             2@                                   �?�q�q�?             "@        ������������������������       �                      @                                   Z@؇���X�?             @                                   V@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@                                  �`@�z�G��?             $@        ������������������������       �                      @                !       
             �?      �?              @        ������������������������       �                      @        "       #                   �b@r�q��?             @        ������������������������       �                     @        $       %                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        '       @                    �?�W���?h            @d@        (       /                   `\@&�a2o��?'            @Q@        )       *                    �?��
ц��?             *@        ������������������������       �                     @        +       ,                   �k@�z�G��?             $@        ������������������������       �                     @        -       .                   �b@      �?             @        ������������������������       �                     @        ������������������������       �                     @        0       9                    �?�>4և��?             L@       1       8                    �?�7��?            �C@       2       3                    �?��S�ۿ?             >@        ������������������������       �                     @        4       7       	          @33�?�8��8��?             8@       5       6                    @M@�����?             5@       ������������������������       �                     3@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        :       ;                    h@��.k���?	             1@        ������������������������       �                     @        <       ?                   @`@�	j*D�?             *@        =       >                   �q@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        A       B                   `a@�L��ȕ?A            @W@       ������������������������       �        -            �P@        C       D                    �N@ ��WV�?             :@       ������������������������       �                     9@        ������������������������       �                     �?        F       G                   @^@DX�\��?*            �Q@        ������������������������       �        
             3@        H       I                   �U@��WV��?              J@        ������������������������       �                     ,@        J       K       
             �?�I�w�"�?             C@        ������������������������       �                     @        L       M                   xs@`Jj��?             ?@       ������������������������       �                     <@        N       O       	          @33�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        Q       j                   �d@�B�gO|�?�            �u@        R       g                    �Q@�ʈD��?8            �U@       S       \                    �?xdQ�m��?4            @T@        T       W       
             �?      �?             8@        U       V                   @_@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        X       Y       	          033@�}�+r��?             3@       ������������������������       �        	             0@        Z       [                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ]       b                    c@���U�?&            �L@       ^       _       
             �?p���?!             I@       ������������������������       �                    �F@        `       a                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        c       d       
             �?؇���X�?             @       ������������������������       �                     @        e       f                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        h       i       	          ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        k       �                   �a@&[i`��?�            Pp@       l       s                    �?(N:!���?h            �e@        m       r                    �?����X�?             <@       n       o       	          ����?r�q��?             8@        ������������������������       �                     @        p       q                   @X@���N8�?
             5@        ������������������������       �                     �?        ������������������������       �        	             4@        ������������������������       �                     @        t       �                    �R@Hm_!'1�?[            `b@       u       �                    �?�'g�2�?Y            �a@       v              
             �?`J����?N            �^@       w       ~                   ``@ _�@�Y�?K             ]@        x       }                    \@ �#�Ѵ�?            �E@        y       z       	          033�?�<ݚ�?             "@        ������������������������       �                     �?        {       |       	          ���@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     A@        ������������������������       �        .            @R@        �       �                   �s@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   pg@      �?             4@        ������������������������       �                     �?        �       �                    Y@���y4F�?
             3@        ������������������������       �                      @        �       �                   �s@�t����?	             1@       �       �                   �`@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �]@h�|�`�?6            �U@        �       �                   �k@d}h���?             ,@        ������������������������       �                      @        �       �                   �Z@      �?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?*O���?.             R@        �       �                    �?�����H�?             B@        ������������������������       �                     3@        �       �                   0m@������?             1@        ������������������������       �                      @        �       �                    @J@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �C@b�2�tk�?             B@        ������������������������       �                     @        �       �                   �j@     ��?             @@        �       �                   i@X�<ݚ�?             "@       �       �                    @M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @N@��<b���?             7@       �       �                   hq@      �?             0@       ������������������������       �        	             (@        �       �                    �L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?և���X�?             @        ������������������������       �                      @        �       �                   �b@z�G�z�?             @        �       �                   m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  ��X�5�?��S�$e�?�5eMYS�?֔5eMY�?�@T:�g�?���7a�?�u�{���?�E(B�?      �?        ��Moz��?Y�B��?      �?        ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?      �?              �?      �?      �?      �?              �?      �?              �?        ��	���?����L�?;�;��?;�;��?�־a�?A��)A�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?ffffff�?333333�?              �?      �?      �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �tk~X��?~X�<ݺ?��Q�g��?ہ�v`��?�;�;�?�؉�؉�?              �?ffffff�?333333�?      �?              �?      �?      �?                      �?�$I�$I�?�m۶m��?��[��[�?�A�A�?�������?�?      �?        UUUUUU�?UUUUUU�?=��<���?�a�a�?      �?                      �?      �?              �?        �������?�?              �?vb'vb'�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        ��~���?X`��?      �?        O��N���?;�;��?      �?                      �?�D+l$�?�]�����?              �?��؉���?��N��N�?              �?����k�?�5��P�?              �?���{��?�B!��?      �?        UUUUUU�?UUUUUU�?              �?      �?        re��?d���y�?�}A_з?A_���?X�<ݚ�?�5?,R�?      �?      �?�������?333333�?              �?      �?        (�����?�5��P�?              �?UUUUUU�?UUUUUU�?              �?      �?        p�}��?	�#����?{�G�z�?\���(\�?              �?�������?�������?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        333333�?�������?              �?      �?        �C��:��?/�I��?�A�A�?|�W|�W�?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?        �a�a�?��y��y�?      �?                      �?      �?        9/���?Y�Cc�?�^���?$T�ik��?�h
���?�~Y���?�{a���?#,�4�r�?�}A_Ч?�/����?�q�q�?9��8���?      �?              �?      �?              �?      �?                      �?              �?�$I�$I�?�m۶m��?              �?      �?              �?      �?      �?        (������?6��P^C�?      �?        �?<<<<<<�?      �?      �?              �?      �?              �?              �?      �?              �?      �?        ⎸#��?��#�;�?I�$I�$�?۶m۶m�?      �?              �?      �?              �?333333�?�������?              �?      �?        �q�q�?�q�q�?�q�q�?�q�q�?              �?�?xxxxxx�?              �?�q�q�?r�q��?              �?      �?        �8��8��?9��8���?              �?      �?      �?�q�q�?r�q��?�������?�������?      �?                      �?              �?��,d!�?��Moz��?      �?      �?      �?              �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��nhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKǅ�h��B�1         �       
             �?"�\�&U�?�           ��@                                 0b@,%�L���?            {@                                  �c@��Y��]�?I            �^@                                 `f@ ����?F            �]@                                 �]@�6H�Z�?D            @]@        ������������������������       �        "            @P@               
                   @^@ pƵHP�?"             J@               	                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �F@                                    O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?               7                    �?þ�%��?�            ps@               ,                   �b@h�����?)             L@              +                    �P@:ɨ��?            �@@                                  �?r֛w���?             ?@                      	          ����?      �?	             $@        ������������������������       �                     @                      	          033�?����X�?             @                                  @      �?             @                     	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               &       	          033�?؇���X�?             5@               %                    �?      �?	             0@       !       $                   �^@@4և���?             ,@        "       #       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        '       *       	             @���Q��?             @        (       )                     I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        -       6                   �b@�LQ�1	�?             7@       .       5       	          ���@�t����?             1@       /       4       	          ����?      �?             0@        0       1                    �J@      �?             @        ������������������������       �                      @        2       3                   @a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             (@        ������������������������       �                     �?        ������������������������       �                     @        8       a                    �?Rq�����?�            �o@       9       J       	          ����?x�f�'�?q            `f@        :       ;       	            �?�MWl��?#            �L@        ������������������������       �                     9@        <       C                    �?     ��?             @@        =       >                    @H@r�q��?             (@        ������������������������       �                     �?        ?       @       	             �?�C��2(�?             &@       ������������������������       �                     @        A       B                    �M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        D       I                   �[@R���Q�?             4@        E       F                    �J@      �?             @        ������������������������       �                      @        G       H                   �Z@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        K       L                   �Z@ �p���?N            �^@        ������������������������       �                      @        M       `                   �e@�(\����?M             ^@       N       _       	          ��� @ ����?L            �]@       O       P       	          `ff�?�J�T�?-            �Q@        ������������������������       �                     .@        Q       R       
             �?h�����?%             L@        ������������������������       �                     @        S       Z       	          ����?�&=�w��?$            �J@        T       U                    �?$�q-�?             *@        ������������������������       �                     �?        V       Y                    @F@�8��8��?             (@        W       X                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             $@        [       \                    q@�(\����?             D@       ������������������������       �                     ;@        ]       ^                   8q@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     H@        ������������������������       �                     �?        b       y                   �d@���=A�?2             S@       c       f       
             �?�w��@�?*            �O@        d       e                   �^@      �?              @        ������������������������       �                      @        ������������������������       �                     @        g       x       	          ����?"pc�
�?&            �K@       h       q       	          ����?�t����?             A@       i       l                   p@r�q��?             8@       j       k                   �i@�X�<ݺ?             2@        ������������������������       �                     �?        ������������������������       �        
             1@        m       p                   �b@      �?             @        n       o                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        r       u       	          ����?���Q��?	             $@       s       t                   �[@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        v       w                   �^@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        z                          �`@�	j*D�?             *@       {       |                    �F@      �?              @       ������������������������       �                     @        }       ~                   `]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    r@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    P@�\m����?�            �r@        �       �       	          ����?ܷ��?��?             =@        �       �                   �Y@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���N8�?             5@        ������������������������       �                      @        �       �                    �?$�q-�?             *@       ������������������������       �                     &@        �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��Lu-��?�            �p@       �       �       	          033@0 �����?�            @n@       �       �                     L@X�aC�U�?�            �m@       �       �       	          pff�?��8����?             h@       �       �                    �?�����?r            �e@        �       �                    �I@�Ń��̧?             E@       ������������������������       �                     B@        �       �                    @J@r�q��?             @        �       �                   0c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        Y            ``@        �       �                   �c@���y4F�?             3@        ������������������������       �                     �?        �       �                   �_@r�q��?             2@        �       �                   �g@և���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �Y@t/*�?             �G@        ������������������������       �                     �?        �       �                   �b@*
;&���?             G@       ������������������������       �                     6@        �       �                    a@�q�q�?             8@        �       �                    @�q�q�?             @       �       �                   Pe@���Q��?             @       �       �                    �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �d@r�q��?
             2@       �       �       	             �?և���X�?             @       �       �                    �M@���Q��?             @        �       �                    �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        �       �                    �?l��[B��?             =@        ������������������������       �                     @        �       �                   �d@�X����?             6@       �       �       	          ����?�t����?             1@        �       �                   �a@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�Bp  ��j��`�?:�J;�O�?��S���?V�����?������?8��18�?�5�5�?�Qv�Qv�?���?�������?              �?;�;��?'vb'vb�?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?      �?      �?                      �?      �?      �?              �?      �?        �����?D;�� �?%I�$I��?n۶m۶�?e�M6�d�?N6�d�M�?�B!��?���{��?      �?      �?      �?        �$I�$I�?�m۶m��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�$I�$I�?۶m۶m�?      �?      �?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        Nozӛ��?d!Y�B�?<<<<<<�?�?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?                      �?              �?�������?�������?���X6��?(��49��?�YLg1�?:��,���?              �?      �?      �?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?        �������?�������?      �?                      �?333333�?333333�?      �?      �?              �?      �?      �?              �?      �?                      �?������?�>�%C��?      �?        �������?333333�?�5�5�?�Qv�Qv�?��V؜?(�K=�?              �?�$I�$I�?�m۶m��?              �?�x+�R�?tHM0���?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�������?333333�?              �?;�;��?�؉�؉�?      �?                      �?              �?      �?        �P^Cy�?��P^Cy�?AA�?�}��}��?      �?      �?              �?      �?        F]t�E�?/�袋.�?�������?�������?UUUUUU�?�������?�q�q�?��8��8�?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?333333�?�������?�������?�������?              �?      �?        �������?333333�?      �?                      �?              �?vb'vb'�?;�;��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?              �?      �?        �Q����?R���Q�?a���{�?��=���?      �?      �?              �?�������?333333�?      �?              �?      �?              �?      �?        �a�a�?��y��y�?              �?;�;��?�؉�؉�?              �?      �?      �?              �?      �?        �X>b�V�?�9�H�?n,�Ra��?���k��?���hB�?Tn�wp٫?�����*�?�������?&>��?���"�w?��<��<�?�a�a�?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?              �?        6��P^C�?(������?              �?�������?UUUUUU�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?              �?        �;����?W�+���?              �?���,d!�?8��Moz�?      �?        �������?�������?UUUUUU�?UUUUUU�?�������?333333�?      �?      �?              �?      �?              �?                      �?�������?UUUUUU�?�$I�$I�?۶m۶m�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?                      �?GX�i���?���=��?      �?        ]t�E]�?�E]t��?�?<<<<<<�?�$I�$I�?�m۶m��?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJXk�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK߅�h��B�7         �                    �?�����?�           ��@              s                   �u@��5Е��?�             y@              h                   �c@\n(�l��?�            @x@              /       
             �?�֞�%��?�            �t@                                  Z@�d2 Λ�?�            �i@        ������������������������       �                     C@               .                    �?�/ C-��?t            �d@                                  �?6�`��V�?V             _@        	                          @c@D�n�3�?             3@       
                           �?     ��?             0@        ������������������������       �                     @                                   �G@      �?             $@        ������������������������       �                     @                                  �s@����X�?             @                                  �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               -       	          ����?(N:!���?I            @Z@              ,                   �b@$gv&��?)            �M@              +                   pb@������?            �F@              "                   `_@d}h���?             E@                                  �O@�����H�?             ;@                                 �k@�}�+r��?             3@       ������������������������       �                     ,@                                   �K@z�G�z�?             @                                  �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                !                     P@      �?              @        ������������������������       �                      @        ������������������������       �                     @        #       (                    `@���Q��?
             .@        $       %                    �E@r�q��?             @        ������������������������       �                     @        &       '                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        )       *                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        ������������������������       �                      G@        ������������������������       �                     E@        0       G                   �f@���@M^�?C             _@        1       F                   �b@     ��?             H@       2       E                    �?�	j*D�?            �C@       3       B                   �d@
;&����?             7@       4       5                   �\@ҳ�wY;�?	             1@        ������������������������       �                     @        6       7                   �X@      �?             (@        ������������������������       �                      @        8       A                   �b@���Q��?             $@       9       @                   �`@      �?              @       :       ;                   `\@؇���X�?             @        ������������������������       �                     @        <       ?                    �?      �?             @       =       >       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        C       D                   �e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        ������������������������       �                     "@        H       g       	          ����?�w�"w��?)             S@       I       R                   �a@<ݚ�?'             R@        J       O                     P@��a�n`�?             ?@       K       L                    �K@ 7���B�?             ;@       ������������������������       �                     2@        M       N                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        P       Q                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        S       X                   @c@#z�i��?            �D@        T       U       	          ����?�����H�?             "@        ������������������������       �                     @        V       W                   �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Y       \                    �?     ��?             @@        Z       [                    �L@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ]       ^                   �i@      �?             8@        ������������������������       �                     �?        _       `                   �l@���}<S�?             7@        ������������������������       �                     $@        a       f       	          @33�?8�Z$���?             *@       b       c                   �c@z�G�z�?             $@        ������������������������       �                     @        d       e                   `p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        i       j                    �O@(;L]n�?"             N@       ������������������������       �                     I@        k       r                    �?z�G�z�?             $@       l       q                    �Q@�q�q�?             @       m       n                    �?z�G�z�?             @        ������������������������       �                     �?        o       p                   Hq@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        t       {                   �`@����X�?             ,@        u       v                    @J@      �?             @        ������������������������       �                      @        w       x       
             �?      �?             @        ������������������������       �                      @        y       z                     O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        |       �                    �?      �?              @       }       �       
             �?؇���X�?             @        ~                           b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �K@���Fi�?�            �t@       �       �                    �?\�����?�            @j@       �       �       
             �?�[|x��?{            �g@        �       �                     B@����e��?            �@@        ������������������������       �                     @        �       �                    ]@8^s]e�?             =@        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?"pc�
�?             6@       �       �       	          ����?�IєX�?             1@        ������������������������       �                     $@        �       �                   @l@؇���X�?             @        ������������������������       �                     @        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@���Q��?             @       �       �                   pj@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �I@�(�Tw�?d            �c@       ������������������������       �        F            �Z@        �       �                    �?`2U0*��?             I@       ������������������������       �                     ?@        �       �                   �U@�KM�]�?             3@        ������������������������       �                      @        ������������������������       �                     1@        �       �       	          hff�?�ՙ/�?             5@        �       �       
             �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?      �?	             ,@        ������������������������       �                     @        �       �                    �?�z�G��?             $@        ������������������������       �                     @        �       �                     H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��\j���?M            �^@        �       �                    �?��a�n`�?             ?@        �       �       	          ����?      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �X@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        �       �       
             �?��+�ޯ�?;            �V@       �       �                    @O@���h%��?)            �O@       �       �       
             �?� ��1�?            �D@        �       �                     N@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �r@�MI8d�?            �B@       �       �                    @L@؇���X�?            �A@        �       �                    _@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?$�q-�?             :@       �       �                    @N@�t����?             1@        ������������������������       �                      @        �       �                   0b@�<ݚ�?             "@       �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�eP*L��?             6@       �       �                   pm@����X�?             ,@       �       �       	          ����?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                   �j@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    U@      �?             <@        ������������������������       �                     @        �       �       	          hff @�J�4�?             9@       �       �                    c@���}<S�?             7@       ������������������������       �                     3@        �       �                   �m@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ������?�v
��,�?*g���?�jL�*�?�W?��? tT����?Q��+Q�?W�v%jW�?�����ܼ?dddddd�?              �?"�%��?8�:����?���{��?B!��?l(�����?(������?      �?      �?      �?              �?      �?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?              �?                      �?�A�A�?|�W|�W�?��/���?[4��}�?�?wwwwww�?۶m۶m�?I�$I�$�?�q�q�?�q�q�?(�����?�5��P�?              �?�������?�������?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?�������?333333�?�������?UUUUUU�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?              �?      �?              �?                      �?              �?              �?�s�9��?�c�1��?      �?      �?;�;��?vb'vb'�?Y�B��?�Mozӛ�?�������?�������?      �?              �?      �?              �?333333�?�������?      �?      �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?      �?                      �?      �?                      �?              �?UUUUUU�?�������?              �?      �?                      �?      �?        ���k(�?��k(��?�q�q�?��8��8�?�s�9��?�c�1Ƹ?	�%����?h/�����?      �?        �q�q�?�q�q�?              �?      �?              �?      �?      �?                      �?�+Q��?ە�]���?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?      �?              �?ӛ���7�?d!Y�B�?      �?        ;�;��?;�;��?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�?�������?              �?�������?�������?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?              �?      �?              �?                      �?�m۶m��?�$I�$I�?      �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        �C.+J�?��FS���?��~��~�?��	��	�?]�u]�u�?EQEQ�?e�M6�d�?6�d�M6�?              �?|a���?	�=����?�$I�$I�?�m۶m��?      �?                      �?/�袋.�?F]t�E�?�?�?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?      �?      �?              �?      �?              �?        p��o���?�A�A�?      �?        ���Q��?{�G�z�?      �?        �k(���?(�����?              �?      �?        �<��<��?�a�a�?۶m۶m�?�$I�$I�?              �?      �?              �?      �?              �?ffffff�?333333�?      �?              �?      �?      �?                      �?�����?�d����?�c�1��?�s�9��?      �?      �?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �Mozӛ�?d!Y�B�?              �?      �?        ]��\���?R�Q��?EQEQ�?v]�u]��?������?������?      �?      �?      �?                      �?L�Ϻ��?��L���?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?;�;��?�؉�؉�?�?<<<<<<�?              �?�q�q�?9��8���?      �?      �?              �?      �?              �?                      �?      �?      �?      �?                      �?t�E]t�?]t�E�?�m۶m��?�$I�$I�?]t�E�?F]t�E�?              �?      �?                      �?      �?      �?      �?                      �?      �?      �?              �?�z�G��?{�G�z�?ӛ���7�?d!Y�B�?      �?              �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ0��JhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKۅ�h��B�6         d       	          ����?0����?�           ��@                                 �`@�I{A�?�            �x@                                  �W@      �?.             T@        ������������������������       �                     6@                                  �c@д>��C�?#             M@                     
             �?��x_F-�?             �I@                                  �?��?^�k�?            �A@       ������������������������       �                     ;@        	                           �?      �?              @       
              	          ���ٿz�G�z�?             @        ������������������������       �                      @                                   \@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                   �?     ��?             0@                                  �?"pc�
�?             &@                                 �]@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               A                    �K@L�Sg��?�            �s@                                  �A@8��T;��?�            �m@                      
             �?և���X�?             ,@        ������������������������       �                     @        ������������������������       �                      @               0       
             �?�>4և��?�             l@               )                    �?�q�q�?             H@              &       	          833�?�q�q�?             8@               !                   �b@�X�<ݺ?             2@       ������������������������       �        	             ,@        "       #                   l@      �?             @        ������������������������       �                      @        $       %                     I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        '       (                   �p@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        *       +                    @G@      �?             8@       ������������������������       �                     &@        ,       -                   �n@�	j*D�?             *@        ������������������������       �                     @        .       /                   �_@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        1       4                   �e@�C��2(�?p             f@        2       3                    �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        5       @                    `@@ o����?j            �d@       6       7                   �c@ qP��B�?6            �U@       ������������������������       �        #             O@        8       =                   �_@�8��8��?             8@       9       <                    �?���7�?             6@        :       ;                     I@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     2@        >       ?                    @H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        4            �S@        B       G                    _@
j*D>�?0            �S@        C       F                    Z@�E��ӭ�?             2@       D       E       
             �?�q�q�?	             (@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        H       [                   �r@�q�q�?"             N@       I       X                    �?�7����?            �G@       J       K                   �a@>��C��?            �E@        ������������������������       �                     .@        L       W                     O@X�Cc�?             <@       M       V                    b@�\��N��?             3@       N       O       	          @33�?      �?             (@        ������������������������       �                     @        P       Q                   b@      �?             @        ������������������������       �                      @        R       U                   pc@      �?             @       S       T                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        Y       Z                   pc@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        \       ]                    t@��
ц��?             *@        ������������������������       �                     @        ^       c                    �?�q�q�?             "@       _       b                    �?      �?              @        `       a                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        e       �       	          ���@��}� �?�             u@       f       �                   P`@�s�>���?�            �p@       g       r                   �\@���Ȓ��?n            `d@        h       i                   �R@���Q��?             4@        ������������������������       �                     @        j       q                   �p@�n_Y�K�?             *@       k       p       	          ����?z�G�z�?             $@       l       m                    �?�����H�?             "@       ������������������������       �                     @        n       o                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        s       �                    f@@2����?`            �a@       t       �                   �]@���۟�?]            `a@       u       x                   �Q@ qP��B�?8            �U@        v       w                   �l@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        y       �                    �?����ȫ�?6            �T@       z       {                    t@�h����?&             L@       ������������������������       �        #            �I@        |                           @M@z�G�z�?             @       }       ~       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        �       �                    ^@f1r��g�?%            �J@        �       �                   �s@�	j*D�?             *@       �       �                    �?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        �       �                    �D@ףp=
�?             D@        �       �                    b@����X�?             @       ������������������������       �                     @        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�FVQ&�?            �@@       ������������������������       �                     :@        �       �       
             �?����X�?             @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @       �       �                    �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          pff�?�ɭ�BR�?H            �Y@        �       �                    �?�[�IJ�?             �G@       �       �       
             �?�q�q�?             8@        ������������������������       �                      @        �       �       	          033�?�GN�z�?             6@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                    �K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?      �?             0@        �       �                   �f@�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �n@�LQ�1	�?             7@       �       �                    �?      �?             (@       �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �       	          033�?z�G�z�?             @        ������������������������       �                     �?        �       �                   �m@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �?Dc}h��?(             L@        ������������������������       �        
             ,@        �       �                   0o@�D����?             E@       �       �                     Q@�������?             >@       �       �                    �F@V�a�� �?             =@        ������������������������       �                     @        �       �                   @e@��+7��?             7@       �       �                     J@��s����?             5@        �       �                   �j@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?�����H�?             2@        �       �       	          `ff�?����X�?             @        ������������������������       �                     @        �       �                   pb@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@r�q��?	             (@       �       �                    a@�C��2(�?             &@       ������������������������       �                     @        �       �                   �a@      �?             @       �       �                   b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�k~X��?+             R@       ������������������������       �                      I@        �       �                   �_@���7�?             6@        �       �                     K@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ���^L�?���Y�?[�R�֯�?K�Z�R��?      �?      �?              �?|a���?a���{�?�?�������?�A�A�?_�_��?              �?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?/�袋.�?F]t�E�?      �?      �?      �?                      �?      �?                      �?              �?ӑ=Q��?��	�Z�?+t+t�?T/�S/��?�$I�$I�?۶m۶m�?              �?      �?        %I�$I��?n۶m۶�?�������?�������?�������?UUUUUU�?�q�q�?��8��8�?              �?      �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?        ;�;��?vb'vb'�?              �?�$I�$I�?۶m۶m�?      �?                      �?t�E]t�?t�E]t�?]t�E�?F]t�E�?              �?      �?        �?�����?�0�ӈ?��}A�?�}A_З?      �?        UUUUUU�?UUUUUU�?�.�袋�?F]t�E�?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?        b'vb'v�?;�;��?r�q��?�q�q�?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?]AL� &�?G}g����?$�;��?qG�w��?      �?        %I�$I��?�m۶m��?�5��P�?y�5���?      �?      �?      �?              �?      �?              �?      �?      �?      �?      �?              �?      �?              �?                      �?      �?              �?      �?              �?      �?        �؉�؉�?�;�;�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?              �?                      �?�n_Y�K�?[$��m�?0{���?�g	�?�E:i�?�\w���?�������?333333�?              �?;�;��?ى�؉��?�������?�������?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?-)D�{�?�7�P�?����j�?��a����?�}A_З?��}A�?      �?      �?              �?      �?        ������?������?�$I�$I�?۶m۶m�?              �?�������?�������?      �?      �?      �?                      �?              �?              �?�x+�R�?�!5�x+�?;�;��?vb'vb'�?F]t�E�?/�袋.�?              �?      �?              �?        �������?�������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?|���?>����?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?��">�T�?ch���V�?m�w6�;�?���
b�?�������?�������?              �?�袋.��?]t�E�?      �?      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?        Y�B��?��Moz��?      �?      �?�������?�������?              �?�������?�������?              �?      �?      �?              �?      �?              �?                      �?�$I�$I�?۶m۶m�?      �?        �0�0�?z��y���?�������?�������?��{a�?a���{�?      �?        zӛ����?Y�B��?z��y���?�a�a�?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?UUUUUU�?�������?F]t�E�?]t�E�?              �?      �?      �?      �?      �?              �?      �?                      �?      �?        �q�q�?�8��8��?              �?F]t�E�?�.�袋�?      �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJڡWhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKɅ�h��B@2         j       	          ����?4�5����?�           ��@              /       
             �?�q�q�?�            @w@                      	          833�?      �?Z            �`@              	                    �?�_�s���?G            @Y@                                  �?��v$���?+            �N@                                   �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        %             K@        
                           @L@�z�G��?             D@                                 @b@X�<ݚ�?             ;@                                 �^@z�G�z�?
             .@                                 `]@�q�q�?             "@                                  �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                  �`@      �?             (@                                  �?      �?             @                                  �?���Q��?             @        ������������������������       �                      @                                  `]@�q�q�?             @        ������������������������       �                     �?                                  �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             *@                                   `_@f���M�?             ?@        ������������������������       �                     @        !       "                    �?������?             ;@        ������������������������       �                     &@        #       .                    �?     ��?             0@       $       %                    �?X�Cc�?	             ,@        ������������������������       �                     @        &       '                     J@X�<ݚ�?             "@        ������������������������       �                     @        (       )                   �_@�q�q�?             @        ������������������������       �                      @        *       +                   �b@      �?             @        ������������������������       �                     �?        ,       -                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        0       Q                    �L@8��8���?�             n@       1       :                    �?��S�ۿ?}            `h@        2       7                    �E@V�a�� �?             =@        3       6                    �?      �?              @       4       5                     C@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        8       9                   �b@���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?        ;       L       	          833�?x�}���?l            �d@       <       ?                   @E@p���?a            �b@        =       >                    �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        @       A                   �l@`׀�:M�?_            �b@       ������������������������       �        0            @S@        B       I                    �?�J�T�?/            �Q@       C       H                    \@ ��ʻ��?-             Q@        D       G                    �?z�G�z�?             @        E       F                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        (            �O@        J       K                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        M       N                    �E@      �?             0@        ������������������������       �                     @        O       P                   �Z@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        R       i       	          ����?������?             �F@       S       d                    �?d}h���?             E@        T       U                   �Y@�q�q�?             8@        ������������������������       �                     �?        V       c       	          ����?8����?             7@       W       b                   Pd@j���� �?	             1@       X       Y                    �?�q�q�?             (@        ������������������������       �                     @        Z       [                    �?����X�?             @        ������������������������       �                     �?        \       a       	          ����?�q�q�?             @       ]       ^                   �_@z�G�z�?             @        ������������������������       �                      @        _       `                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        e       f                    �O@�X�<ݺ?             2@       ������������������������       �                     (@        g       h                    s@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        k       �                    �?������?�            �v@       l       �       
             �?Pe6�p�?�            �p@       m       �                    c@���,�g�?�            `l@       n       w                    j@T�y���?|            `j@        o       t                   i@v���a�?*            @R@       p       q                   Pe@`Jj��?%             O@       ������������������������       �                    �G@        r       s                   �e@������?	             .@        ������������������������       �                     @        ������������������������       �                     &@        u       v                   �`@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        x       �                    `R@��.N"Ҭ?R            @a@       y       �       	          ����?`Y����?Q             a@        z       {       
             �?R���Q�?             4@        ������������������������       �                     �?        |       }                   8r@�KM�]�?             3@       ������������������������       �        
             (@        ~       �                    �?����X�?             @              �                   �_@r�q��?             @        ������������������������       �                     @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        B            @]@        ������������������������       �                     �?        �       �                    �?     ��?             0@       �       �                    @O@      �?              @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?^H���+�?            �B@        �       �                    �J@d}h���?             ,@        �       �                   0a@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �`@���}<S�?             7@       �       �                    �?8�Z$���?             *@        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                     Q@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �       
             �?�`���??            �X@       �       �                    �?���Q��?.            �Q@        �       �                    �M@$�q-�?	             *@       ������������������������       �                     $@        �       �                    @P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @��h!��?%            �L@       �       �       	          `ff�?~���L0�?            �H@       �       �                   �l@      �?             :@       �       �                   �Z@�q�q�?
             2@        ������������������������       �                     @        �       �                   �`@z�G�z�?             .@       ������������������������       �                     "@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                   �r@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���}<S�?             7@        �       �                   @_@      �?             @        ������������������������       �                     �?        �       �                   0b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        �       �                    �?      �?              @       �       �                    @L@r�q��?             @        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	          ���@d}h���?             <@       �       �       	          ����?H%u��?             9@       �       �                    �L@���!pc�?	             &@       ������������������������       �                     @        �       �                   n@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�   Np	�?���Gw{�?UUUUUU�?UUUUUU�?      �?      �?Q`ҩy�?��g����?;ڼOqɐ?.�u�y�?�$I�$I�?۶m۶m�?      �?                      �?              �?333333�?ffffff�?�q�q�?r�q��?�������?�������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?      �?                      �?      �?      �?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?                      �?��RJ)��?��Zk���?              �?B{	�%��?{	�%���?      �?              �?      �?%I�$I��?�m۶m��?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?�������?�?��{a�?a���{�?      �?      �?      �?      �?      �?                      �?              �?��y��y�?�a�a�?      �?                      �?�(፦�?4u~�!��?\���(\�?{�G�z�?      �?      �?      �?                      �?��L��?к����?      �?        (�K=�?��V؜?�������?�?�������?�������?      �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?�؉�؉�?;�;��?              �?      �?        wwwwww�?�?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?              �?d!Y�B�?8��Moz�?�������?ZZZZZZ�?�������?�������?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        ��8��8�?�q�q�?      �?        �������?UUUUUU�?      �?                      �?              �?(��$�?�J�v|�?���>��?�|���?*���ϸ?�*����?�&��2�?&�k]���?�4iҤI�?ٲe˖-�?�B!��?���{��?              �?�?wwwwww�?      �?                      �?]t�E]�?F]t�E�?      �?                      �?ہ�v`��?�3J���?�d�*al�?�,���L�?333333�?333333�?      �?        (�����?�k(���?              �?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?                      �?      �?              �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?              �?      �?        �g�`�|�?L�Ϻ��?I�$I�$�?۶m۶m�?�������?333333�?              �?      �?              �?        d!Y�B�?ӛ���7�?;�;��?;�;��?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?              �?              �?����S�?և���X�?�������?333333�?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        p�}��?Hp�}�?������?����>4�?      �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?              �?      �?              �?      �?              �?      �?        d!Y�B�?ӛ���7�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?I�$I�$�?۶m۶m�?)\���(�?���Q��?F]t�E�?t�E]t�?      �?              �?      �?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:d�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         h       	             �?6�L����?�           ��@              7                    �?p9W��S�?�            �w@                      
             �?�ƥ���?\            �a@                                   �O@     ��?+             P@                                  �?4��?�?$             J@                                   �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        	                           �? qP��B�?            �E@        
                          �c@�X�<ݺ?             2@       ������������������������       �        
             (@                                   �?r�q��?             @                                 �o@      �?             @                                  pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     9@                                  �`@�q�q�?             (@                                  �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               (                   �b@�2��?1            �S@              '       	          ����?�q�q�?             H@              "                    P@�����?             E@               !       	          ����?      �?             @                                  �?      �?             @        ������������������������       �                      @                                   e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        #       &                    �?������?             B@        $       %                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     <@        ������������������������       �                     @        )       2                   @d@`՟�G��?             ?@        *       -                    �?     ��?             0@        +       ,                    s@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        .       /                   �`@�C��2(�?	             &@       ������������������������       �                     "@        0       1                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       6                    �?��S�ۿ?             .@        4       5                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        8       M                    �K@0>�Xu�?�            �m@       9       @                    ]@ �ղ?n            �f@        :       ?                    �?�KM�]�?             C@       ;       <                   �o@�L���?            �B@       ������������������������       �                     :@        =       >                   �p@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        A       B                    @E@@��t��?W             b@        ������������������������       �                      L@        C       H                   `a@X;��?7            @V@       D       G                    �E@ ��ʻ��?'             Q@        E       F                    @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        "             N@        I       J                    �?�����?             5@       ������������������������       �                     ,@        K       L       	          ����?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        N       U                    �?      �?$             K@        O       T                   �c@z�G�z�?             $@       P       Q       
             �?���Q��?             @        ������������������������       �                     �?        R       S                   `r@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        V       c                   �a@~�4_�g�?             F@       W       \                   P`@      �?             @@        X       [                   �_@ףp=
�?             $@        Y       Z       
             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ]       b       
             �?�X����?             6@       ^       _                     Q@      �?             0@       ������������������������       �                     *@        `       a                   pm@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        d       g                    �?�8��8��?             (@        e       f                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        i       �                    �?��mo*�?�             v@        j                          �j@�1�����?S            �`@        k       p                    �?Jm_!'1�?             �H@        l       o                    �P@      �?             $@       m       n                     L@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        q       v                   @[@��-�=��?            �C@        r       s       
             �?�<ݚ�?             "@       ������������������������       �                     @        t       u                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        w       x                    @O@��S�ۿ?             >@       ������������������������       �                     5@        y       z       	          `ff�?�<ݚ�?             "@        ������������������������       �                     �?        {       ~                    @P@      �?              @        |       }                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?t���D�?3            �U@        �       �       
             �?���!pc�?             6@       �       �                   0p@և���X�?             ,@        �       �                   0l@؇���X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          033�?����X�?             @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   @q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �p@     8�?!             P@       �       �                   d@<=�,S��?            �A@       �       �                     P@�㙢�c�?             7@       �       �                   pn@�����?             5@        �       �                    �N@����X�?             @       �       �                    a@r�q��?             @        ������������������������       �                      @        �       �                   �l@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                      @        �       �                   �\@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        �       �       	          ����?д>��C�?             =@       ������������������������       �                     4@        �       �                   �a@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?X��*"�?�            `k@       �       �                   �s@*~k���?f            �b@       �       �                    �?�θV�?]            @a@       �       �                    �F@ ,��-�?P            �]@        �       �                    b@�θ�?	             *@       �       �                   �Z@�C��2(�?             &@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �       �                   Xp@���N8�?G            @Z@       �       �       	          033@@4և���?3            �Q@       �       �       	          033�? 7���B�?(             K@        ������������������������       �                     .@        �       �                    @L@�7��?            �C@        ������������������������       �                     1@        �       �                   `_@�C��2(�?             6@        ������������������������       �                     &@        �       �                   pi@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                   p@     ��?             0@       ������������������������       �        	             &@        �       �                     M@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �A@        �       �                   `_@�z�G��?             4@        ������������������������       �                     &@        �       �                    �?�q�q�?             "@        ������������������������       �                      @        �       �                   p@և���X�?             @       �       �                   �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�	j*D�?	             *@        ������������������������       �                     �?        �       �                    �L@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        �       �                    �R@�IєX�?)             Q@       �       �       	          ����? ����?(            @P@        �       �                   �a@�IєX�?             1@       ������������������������       �                     (@        �       �                   �m@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     H@        ������������������������       �                     @        �t�b��      h�h)h,K ��h.��R�(KK�KK��hb�Bp  6�;����?e���?�k(����?l(�����?$T�ik��?�U0K��?      �?      �?ى�؉��?�N��N��?�q�q�?r�q��?      �?                      �?�}A_З?��}A�?�q�q�?��8��8�?              �?UUUUUU�?�������?      �?      �?      �?      �?      �?                      �?              �?              �?              �?�������?�������?      �?      �?      �?                      �?              �?���JG�?�&��jq�?UUUUUU�?�������?=��<���?�a�a�?      �?      �?      �?      �?      �?              �?      �?      �?                      �?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?�1�c��?�s�9��?      �?      �?�������?333333�?      �?                      �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?�������?�?�������?UUUUUU�?              �?      �?              �?        |!E��h�?z���\�?�/���?��ݮ��?�k(���?(�����?}���g�?L�Ϻ��?      �?        F]t�E�?t�E]t�?              �?      �?                      �?*h���V�?��RA�/�?      �?        �u�{���?�E(B�?�������?�?      �?      �?      �?                      �?      �?        =��<���?�a�a�?      �?        �m۶m��?�$I�$I�?      �?                      �?      �?      �?�������?�������?333333�?�������?              �?      �?      �?      �?                      �?      �?        ��.���?/�袋.�?      �?      �?�������?�������?      �?      �?              �?      �?                      �?]t�E]�?�E]t��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?        W'u_�?�<�"h�?Hֹ�d�?����M�?������?����X�?      �?      �?�$I�$I�?�m۶m��?      �?                      �?      �?        �A�A�?}˷|˷�?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�������?              �?�q�q�?9��8���?      �?              �?      �?      �?      �?              �?      �?                      �?�;⎸�?$�;��?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        �$I�$I�?�m۶m��?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?             ��?      �?X|�W|��?�A�A�?d!Y�B�?�7��Mo�?�a�a�?=��<���?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?                      �?      �?              �?      �?              �?      �?        a���{�?|a���?      �?        �q�q�?r�q��?              �?      �?        x��m���?��C2��?�z=��?��^x/�?�Q�g���?̵s���?'u_[�?[4���?�؉�؉�?ى�؉��?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?      �?        �a�a�?��y��y�?�$I�$I�?n۶m۶�?h/�����?	�%����?              �?�A�A�?��[��[�?              �?F]t�E�?]t�E�?              �?F]t�E�?/�袋.�?      �?                      �?      �?      �?              �?333333�?�������?      �?                      �?              �?333333�?ffffff�?              �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?        ;�;��?vb'vb'�?      �?              �?      �?              �?      �?        �?�? �����? �����?�?�?              �?�������?�������?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�I]fhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�/         �       
             �?������?�           ��@              I                    �?@���^��?           �y@                      
             �?��Y���?e            �c@               	                   �c@������?
             1@                                  �?$�q-�?             *@       ������������������������       �                     "@                                  �X@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        
              	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @               8                    a@:9��z�?[            �a@                                 �R@*u�$��?:            �V@                                   �?���N8�?             5@       ������������������������       �        
             .@                                   @r�q��?             @                                  �K@z�G�z�?             @        ������������������������       �                     @                                  �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                   g@��
P��?+            �Q@        ������������������������       �                     @               3                    �?     ��?(             P@              $                   �a@~h����?$             L@                                   �?�q�q�?             2@        ������������������������       �                     @                                  Pq@$�q-�?	             *@       ������������������������       �                     $@                !                    �G@�q�q�?             @        ������������������������       �                     �?        "       #                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       (                    �?\�Uo��?             C@        &       '                    �K@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        )       .                    �?� �	��?             9@       *       -                   �n@������?
             .@        +       ,                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        /       0                    �K@�z�G��?             $@        ������������������������       �                     @        1       2                   �l@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        4       5                   pb@      �?              @        ������������������������       �                     @        6       7                   �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        9       :                    �?�:pΈ��?!             I@        ������������������������       �                     9@        ;       B       	          833�? �o_��?             9@        <       =                    �?�q�q�?	             (@        ������������������������       �                     @        >       A                    �G@      �?              @        ?       @                   `a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        C       D       	          ����?8�Z$���?	             *@        ������������������������       �                     @        E       F                    W@      �?              @        ������������������������       �                     �?        G       H                    f@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        J       Y                    �?     \�?�             p@        K       X                    �?`՟�G��?             ?@       L       O                    �?��
ц��?             :@        M       N                   0q@      �?              @       ������������������������       �                     @        ������������������������       �                      @        P       S                   �a@X�<ݚ�?	             2@        Q       R                   Pj@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        T       W                   �`@�<ݚ�?             "@        U       V       	          ��� @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        Z       m                   pa@Х-��ٹ?�             l@       [       j                    `P@ qP��B�?W             `@       \       i                   �[@ ����?P            �]@        ]       d                    �?���}<S�?             7@       ^       _                    �K@P���Q�?             4@       ������������������������       �                     *@        `       a                    Y@؇���X�?             @       ������������������������       �                     @        b       c                   �p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        e       h                    �?�q�q�?             @       f       g       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        A             X@        k       l                    �P@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        n       }                    �?     ��?9             X@       o       r                   g@6uH���?%             O@        p       q                   `U@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        s       |                   �b@ �h�7W�?            �J@       t       {                   �a@���J��?            �I@        u       z                    �?���N8�?             5@       v       y                   �l@@4և���?             ,@        w       x       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     >@        ������������������������       �                      @        ~       �       
             �?�t����?             A@               �                   �b@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @N@h�����?             <@       ������������������������       �        
             3@        �       �       	             �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @c@R���	�?�             t@        �       �       	          ����?:ɨ��?            �@@        �       �                   �Y@�	j*D�?	             *@        ������������������������       �                      @        �       �                    �?"pc�
�?             &@       �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?P���Q�?             4@        �       �                     N@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        �       �                    �?D�� ��?�            �q@        �       �                    �?rEC��a�?1            �S@       �       �                     E@6uH���?&             O@        �       �                   �\@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          hff�?h�����?"             L@       ������������������������       �                     H@        �       �                   �d@      �?              @       ������������������������       �                     @        �       �                   0e@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   `l@@�0�!��?             1@        �       �                    �?և���X�?             @        �       �                   `k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                     L@���%�?x             j@       ������������������������       �        a            �d@        �       �                   `d@,���i�?            �D@       �       �                    �?�X�<ݺ?             B@        ������������������������       �                     *@        �       �                    �L@���}<S�?             7@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   ps@���N8�?             5@       ������������������������       �        
             4@        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �sF�v
�?�\��z�?�bPn��?D�{���?-n����?�Ȟ��t�?xxxxxx�?�?�؉�؉�?;�;��?      �?              �?      �?              �?      �?              �?      �?      �?                      �?P$�Ҽ��?����?Z�Z��?�/��/��?�a�a�?��y��y�?              �?UUUUUU�?�������?�������?�������?              �?      �?      �?      �?                      �?              �?PuPu�?_�_��?      �?              �?      �?%I�$I��?�m۶m��?UUUUUU�?UUUUUU�?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�5��P^�?6��P^C�?�؉�؉�?;�;��?      �?                      �?)\���(�?�Q����?�?wwwwww�?UUUUUU�?UUUUUU�?              �?      �?                      �?ffffff�?333333�?      �?              �?      �?              �?      �?              �?      �?              �?      �?      �?              �?      �?        �Q����?��Q���?              �?�Q����?
ףp=
�?�������?�������?      �?              �?      �?      �?      �?      �?                      �?              �?;�;��?;�;��?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?     ��?�s�9��?�1�c��?�;�;�?�؉�؉�?      �?      �?      �?                      �?�q�q�?r�q��?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?9��8���?      �?      �?      �?                      �?              �?              �?O贁N�?K~��K�?�}A_З?��}A�?�5�5�?�Qv�Qv�?d!Y�B�?ӛ���7�?�������?ffffff�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?�������?�������?      �?                      �?      �?      �?��RJ)��?k���Zk�?�q�q�?9��8���?              �?      �?        "5�x+��?��sHM0�?�?______�?�a�a�?��y��y�?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?      �?        �?<<<<<<�?      �?      �?              �?      �?        �$I�$I�?�m۶m��?              �?�q�q�?�q�q�?      �?                      �?�����L�?�������?e�M6�d�?N6�d�M�?vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?�q�q�?�q�q�?      �?                      �?      �?      �?              �?      �?        �������?ffffff�?�$I�$I�?۶m۶m�?              �?      �?                      �?
kxg�R�?��<�\h�?�0���M�?�=Q���?k���Zk�?��RJ)��?      �?      �?              �?      �?        �m۶m��?�$I�$I�?      �?              �?      �?      �?              �?      �?              �?      �?        �������?ZZZZZZ�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?        �������?333333�?      �?                      �?              �?�;�;�?ى�؉��?      �?        �����?8��18�?��8��8�?�q�q�?      �?        ӛ���7�?d!Y�B�?      �?      �?              �?      �?        ��y��y�?�a�a�?      �?                      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�޵#hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKՅ�h��B@5         �       
             �?��}���?�           ��@              M                    �?�Q�G�%�?           0z@               <                    �?���|���?c            �d@                     	          833�?�F�j��?A            �Z@               
                    �?      �?             B@                                   Z@X�<ݚ�?             "@        ������������������������       �                     @               	                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?PN��T'�?             ;@       ������������������������       �                     1@                                   �?���Q��?             $@                                  �b@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?���Q��?             @        ������������������������       �                      @                                  @_@�q�q�?             @                                 0b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                   �G@X�Cc�?)            �Q@                      	             @�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?               )                   �k@��
ц��?!             J@               (       	          ����?��+7��?             7@              %                   �b@��s����?             5@              $       	          033�?      �?
             0@                #                   �g@؇���X�?             @        !       "                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        &       '                   �V@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        *       3                    �?����"�?             =@       +       0                   Xr@�q�q�?             .@       ,       /                   �o@"pc�
�?             &@        -       .                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        1       2       	          033@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        4       9                   �`@և���X�?             ,@        5       8                    �?r�q��?             @       6       7                    @L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        :       ;       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        =       @                    �?�j��b�?"            �M@        >       ?                    d@      �?             @        ������������������������       �                     @        ������������������������       �                     @        A       D       
             �? �h�7W�?            �J@        B       C       	          pff�?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        E       F                    �?`���i��?             F@        ������������������������       �                     @        G       H       	             �?�?�|�?            �B@       ������������������������       �                     ?@        I       J                   �b@r�q��?             @       ������������������������       �                     @        K       L                    e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        N       �                    @4Jı@�?�            �o@       O       ^                    �?X����?�            `o@        P       ]       	          033�?�q�q�?             >@       Q       \                   �s@�G��l��?             5@       R       Y                   �b@D�n�3�?             3@       S       T                    �L@����X�?             ,@        ������������������������       �                     @        U       X                    a@և���X�?             @        V       W                    `@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        Z       [                     K@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        _       �                    �?`���~�?�            �k@       `       �                    �R@ 7���B�?x            �g@       a       x                   pb@�?�|�?v             g@       b       w                    �L@0{�o��?l            @e@       c       j                    \@�zvܰ?8             V@        d       e                   �m@؇���X�?             @        ������������������������       �                     @        f       g                     E@      �?             @        ������������������������       �                      @        h       i                   p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        k       v       	          ����?F|/ߨ�?2            @T@        l       m       	             �?�>����?             ;@        ������������������������       �                     *@        n       u                    m@؇���X�?
             ,@       o       t                    l@      �?              @       p       s                   P`@؇���X�?             @        q       r                   �j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        "             K@        ������������������������       �        4            �T@        y       z       
             �?�r����?
             .@        ������������������������       �                     @        {       |                    \@"pc�
�?             &@        ������������������������       �                     �?        }       ~                   �`@ףp=
�?             $@        ������������������������       �                     @               �                    �?      �?             @        �       �                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �p@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @Y@     ��?             @@        ������������������������       �                      @        �       �                   �`@(;L]n�?             >@       ������������������������       �                     9@        �       �                    @M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?b�h�d.�?�            �s@       �       �                    �?l-MIڼ�?�            0q@       �       �                    �?X�aC�U�?�            �m@        �       �                   �a@r�����?%            �J@        ������������������������       �                     :@        �       �                   `b@��}*_��?             ;@        ������������������������       �                      @        �       �                   �_@`�Q��?             9@        �       �                   0d@�eP*L��?             &@        �       �                   �c@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �       	             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    s@؇���X�?             ,@       ������������������������       �                     $@        �       �                   �c@      �?             @        ������������������������       �                     �?        �       �                   0w@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?0�z��?�?m            @g@        ������������������������       �        +            �R@        �       �                     L@������?B             \@       ������������������������       �        7            @X@        �       �       	          ����?z�G�z�?             .@       ������������������������       �                     "@        �       �       	          ����?      �?             @       �       �                   a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             B@        ������������������������       �                     @        �       �                    �?�z�G��?             >@       �       �                    ]@      �?             <@        ������������������������       �                     @        �       �       	             �? �o_��?             9@        �       �                    h@��
ц��?	             *@        ������������������������       �                     @        �       �                    @J@�q�q�?             "@        �       �                   �e@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          033�?�8��8��?	             (@       ������������������������       �                      @        �       �                   �^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �U@      �?             D@        ������������������������       �        
             2@        �       �                   �`@�C��2(�?             6@       ������������������������       �        	             &@        �       �                   Pc@"pc�
�?             &@       �       �                    �?      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  q��H��?��>���?��ڞ��?CQI�ʼ�?F]t�E�?]t�E]�?��sHM�?:�&oe�?      �?      �?r�q��?�q�q�?              �?�������?UUUUUU�?              �?      �?        h/�����?&���^B�?              �?�������?333333�?�������?�������?      �?                      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?%I�$I��?�m۶m��?��8��8�?�q�q�?      �?                      �?�;�;�?�؉�؉�?zӛ����?Y�B��?z��y���?�a�a�?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �������?333333�?      �?                      �?              �?�i��F�?	�=����?UUUUUU�?UUUUUU�?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?�������?UUUUUU�?�������?�������?              �?      �?              �?              �?      �?      �?                      �?��/���?�N��?      �?      �?              �?      �?        "5�x+��?��sHM0�?�q�q�?9��8���?      �?                      �?F]t�E�?F]t�E�?              �?к����?*�Y7�"�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?��b�X,�?O���t:�?���e�?�_FA@s�?UUUUUU�?UUUUUU�?��y��y�?1�0��?(������?l(�����?�$I�$I�?�m۶m��?              �?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?�������?�������?      �?                      �?      �?                      �?�*�*�??R�>R��?h/�����?	�%����?к����?*�Y7�"�?�?oooooo�?t�E]t�?颋.���?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?      �?      �?                      �?�����H�?�Hx�5�?h/�����?�Kh/��?              �?�$I�$I�?۶m۶m�?      �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?                      �?              �?              �?�?�������?              �?F]t�E�?/�袋.�?      �?        �������?�������?              �?      �?      �?      �?      �?      �?                      �?              �?      �?      �?              �?      �?              �?      �?      �?        �?�������?              �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?;��:���?_�_��?���+�?�j����?���hB�?Tn�wp٫?Dj��V��?�V�9�&�?      �?        _B{	�%�?B{	�%��?              �?��(\���?{�G�z�?]t�E�?t�E]t�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        |���{�?�B!��?      �?        I�$I�$�?۶m۶m�?      �?        �������?�������?      �?              �?      �?      �?      �?              �?      �?              �?        �������?�������?      �?        333333�?ffffff�?      �?      �?              �?�Q����?
ףp=
�?�؉�؉�?�;�;�?              �?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?      �?              �?]t�E�?F]t�E�?      �?        /�袋.�?F]t�E�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�G�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK݅�h��B@7         �       
             �?���:���?�           ��@              {                   �b@ęI0�?           pz@                     	          833�?б��J��?�            �v@                                   �?�kb97�?0            @S@       ������������������������       �                      K@                                  0a@�㙢�c�?             7@                                  `X@���Q��?             $@        ������������������������       �                     �?        	       
                    T@�q�q�?             "@        ������������������������       �                     @                                  @^@���Q��?             @        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             *@               ^                    �?^�R|���?�            r@              E                   �_@2Tv���?�             n@              6                   Pr@`	�<��?[            �a@              -                   `_@�=|+g��?I            @\@              ,                    �?�NW���?D            �Z@                                  �?$��$�L�?1            �S@                                    H@�θ�?             *@        ������������������������       �                     �?                                  @]@r�q��?             (@       ������������������������       �                     @                                   �N@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @               #                    �?�U�=���?)            �P@              "                    `@@3����?!             K@                !                   �_@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     E@        $       )       	             @�q�q�?             (@       %       (                    �L@�<ݚ�?             "@        &       '                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        *       +                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        .       /                    �?����X�?             @        ������������������������       �                      @        0       1                    �?���Q��?             @        ������������������������       �                     �?        2       3       	          ����?      �?             @        ������������������������       �                     �?        4       5       	          033@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        7       @                   �`@��X��?             <@        8       9                    ]@      �?              @        ������������������������       �                     �?        :       ;                   @s@����X�?             @        ������������������������       �                      @        <       =                   @_@���Q��?             @        ������������������������       �                      @        >       ?                   ``@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        A       D                    �Q@z�G�z�?             4@       B       C       	          ����?�����H�?             2@        ������������������������       �                      @        ������������������������       �        
             0@        ������������������������       �                      @        F       I       	          ����?���F6��?;            �X@        G       H                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        J       W                    �?p�qG�?9             X@       K       V       	             �?(;L]n�?4            �V@        L       U                   �`@�8��8��?             B@        M       N                   @_@d}h���?             ,@        ������������������������       �                     �?        O       P       	          ����?8�Z$���?
             *@        ������������������������       �                     �?        Q       R                   `b@�8��8��?	             (@       ������������������������       �                     $@        S       T                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     K@        X       ]                   0`@�q�q�?             @       Y       Z                   @b@      �?             @        ������������������������       �                     �?        [       \                   @q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        _       n                    �?`�(c�?!            �H@        `       m                    �?      �?             8@       a       b                   `Z@���y4F�?             3@        ������������������������       �                     �?        c       l                    �?r�q��?
             2@       d       e                   0g@�t����?	             1@        ������������������������       �                     �?        f       g                   0b@      �?             0@        ������������������������       �                     "@        h       k                    �?؇���X�?             @        i       j                   Pb@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        o       z       	          `ff�?�J�4�?             9@       p       q                    @M@���y4F�?             3@        ������������������������       �                     @        r       y                   �`@�	j*D�?
             *@       s       x                   �s@"pc�
�?             &@       t       w                   �j@ףp=
�?             $@        u       v                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        |       }                    c@���b���?%            �L@        ������������������������       �                     @        ~       �                    �?z�):���?              I@               �                    �?�z�G��?             4@       �       �                   @a@��S�ۿ?	             .@       ������������������������       �                     *@        �       �                   �t@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �f@*;L]n�?             >@       �       �                    @M@`�Q��?             9@       �       �       	          ����?��s����?             5@       ������������������������       �        	             &@        �       �                   �o@���Q��?             $@        �       �                   �c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    S@4�Q�]�?�            ps@        ������������������������       �                      @        �       �       	          ����?�N�_��?�            Ps@       �       �                    @M@Nި*:�?�            �q@       �       �                    �?io8�?�             m@        �       �                   @\@�S����?             C@        �       �                   g@�q�q�?             (@        ������������������������       �                      @        �       �                    �G@z�G�z�?             $@        �       �                   Pd@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @c@$�q-�?             :@        �       �                   �`@�q�q�?             @       �       �                    @H@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �       	            �?��8�$>�?w            @h@       �       �                    @A@@�E��@�?h            �e@        �       �                   �[@�8��8��?             (@        ������������������������       �                     @        �       �                   Pc@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �o@�dJ�Ҙ?a            `d@       ������������������������       �        C             \@        �       �                    �?`'�J�?            �I@       ������������������������       �                    �H@        ������������������������       �                      @        �       �                   `X@�d�����?             3@        ������������������������       �                     @        �       �                    @L@      �?             0@       �       �                    �?��S�ۿ?             .@        �       �                   0l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     �?        �       �                    `R@ڡR����?            �H@       �       �                    �?�L�lRT�?            �F@        �       �                    V@�t����?             1@        ������������������������       �                     @        �       �                    �?      �?             $@        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   Pc@؇���X�?             <@       ������������������������       �        
             2@        �       �                   ht@���Q��?             $@       �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?X�Cc�?             <@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�GN�z�?             6@       �       �       	          ����?�q�q�?             .@        ������������������������       �                     @        �       �                    n@      �?	             $@       �       �                   `]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �G@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  !��Q��?p��1W-�?�k���?e����?�f�"�?Nx��A��?�cj`?�Y�	qV�?              �?d!Y�B�?�7��Mo�?�������?333333�?      �?        UUUUUU�?UUUUUU�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�W��H��?�@�m�?�������?�������?E�)͋?�?o����?Vzja���?���S+�?�x+�R�?萚`���?�3���?��]-n��?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?              �?�������?333333�?              �?      �?        e�M6�d�?�M6�d��?h/�����?���Kh�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?�m۶m��?              �?�������?333333�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?%I�$I��?n۶m۶�?      �?      �?              �?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�q�q�?�q�q�?      �?                      �?      �?        ogH���?�v�ļ�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?�?�������?UUUUUU�?UUUUUU�?۶m۶m�?I�$I�$�?      �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?4և����?������?      �?      �?6��P^C�?(������?              �?�������?UUUUUU�?<<<<<<�?�?              �?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?                      �?              �?{�G�z�?�z�G��?(������?6��P^C�?              �?;�;��?vb'vb'�?F]t�E�?/�袋.�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?                      �?g1��t�?1��t��?      �?        H�z�G�?q=
ףp�?ffffff�?333333�?�������?�?      �?              �?      �?              �?      �?                      �?�������?""""""�?{�G�z�?��(\���?�a�a�?z��y���?              �?�������?333333�?      �?      �?              �?      �?        UUUUUU�?�������?              �?      �?              �?              �?        ��oH�q�?�4@ޞ9�?              �?:�7i��?��![��?�{8� �?� <n���?|a���?GX�i��?(������?^Cy�5�?UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?      �?        �Q�/��?����?ĦҐs�?E'�卑?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        w��|��?)��I� �?      �?        �������?�?      �?                      �?Cy�5��?y�5���?              �?      �?      �?�������?�?      �?      �?              �?      �?              �?                      �?����S��?����X�?�I��I��?l�l��?�������?�������?              �?      �?      �?              �?�m۶m��?�$I�$I�?333333�?�������?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        333333�?�������?۶m۶m�?�$I�$I�?      �?                      �?              �?              �?�m۶m��?%I�$I��?�������?UUUUUU�?      �?                      �?]t�E�?�袋.��?UUUUUU�?UUUUUU�?              �?      �?      �?�������?�������?              �?      �?        �������?�������?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���JhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@+         j                    �?�$���?�           ��@              3       	          ����?�Ǹ6=�?�            `{@                                  @^@d\@som�?Y            �c@                      
             �?���*�?              N@                                 @[@`Ӹ����?            �F@       ������������������������       �                     ?@                                  �`@؇���X�?             ,@        ������������������������       �                     "@        	       
                    �?���Q��?             @        ������������������������       �                      @                                   @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �]@���Q��?             .@                     	          ����?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @                      
             �?��ga�?9            @X@                                   �?�����?             C@                                   �?���|���?             &@                                 �p@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                      	          433�?�+$�jP�?             ;@       ������������������������       �                     6@        ������������������������       �                     @               *                    �?��mo*�?"            �M@                                  �?8��8���?             H@        ������������������������       �                     @                !                   @E@X�EQ]N�?            �E@        ������������������������       �                      @        "       #                    Z@��p\�?            �D@        ������������������������       �                     �?        $       %                   �b@P���Q�?             D@       ������������������������       �                     4@        &       '                   �j@ףp=
�?	             4@        ������������������������       �                     �?        (       )                   `\@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        +       .                    �?"pc�
�?             &@       ,       -                   �`@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        /       2                   �b@�q�q�?             @       0       1                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        4       K                    _@h?\P��?�            �q@        5       B                   �o@z�G�z�?%            �Q@       6       7       
             �?`2U0*��?             I@        ������������������������       �        	             1@        8       9                   `_@�FVQ&�?            �@@        ������������������������       �        	             2@        :       ?                    �K@�r����?
             .@       ;       >                    Z@$�q-�?             *@        <       =       	          ���@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        @       A                   Pl@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        C       J                   �t@���Q��?	             4@       D       I                    �J@�t����?             1@       E       F                   `^@$�q-�?             *@       ������������������������       �                     $@        G       H       	             @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        L       g                    `R@�!ʉ�?t            `j@       M       `       
             �? ��WV�?r             j@       N       O                   `R@`��Zש?h             h@        ������������������������       �                     �?        P       Q                    @L@@��8��?g             h@        ������������������������       �        1             W@        R       _                   �a@`2U0*��?6             Y@       S       Z                   pa@�8��8��?             H@       T       Y                    �L@��?^�k�?            �A@        U       V                    e@z�G�z�?             @        ������������������������       �                     @        W       X       	          033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@        [       \                    a@�θ�?             *@        ������������������������       �                     @        ]       ^                   �c@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     J@        a       b                    �?z�G�z�?
             .@        ������������������������       �                     @        c       f                   p`@      �?             (@        d       e                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        h       i                   �p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       �       
             �?x�Ӵ�q�?�            �r@        l       �                   0`@�f��`��?B            �[@        m       |                   �r@��P���?            �D@       n       {                     P@��hJ,�?             A@       o       z                    @L@`Jj��?             ?@       p       q                   `]@      �?
             0@        ������������������������       �                     @        r       s                    �?"pc�
�?             &@        ������������������������       �                     �?        t       y                    �?ףp=
�?             $@        u       v                    �?r�q��?             @        ������������������������       �                     @        w       x                   �Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     @        }       ~                    Z@և���X�?             @        ������������������������       �                      @               �                    @M@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �e@�z�G��?*            �Q@       �       �                    �G@      �?$             N@        ������������������������       �        
             3@        �       �                    �?��]�T��?            �D@        ������������������������       �                     "@        �       �                   �c@     ��?             @@       �       �       	          `ff�?
j*D>�?             :@       �       �                    �?D�n�3�?             3@        �       �       	          ����?      �?              @        ������������������������       �                     @        �       �       	            �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �j@���|���?	             &@        ������������������������       �                     @        �       �                   �a@      �?              @        ������������������������       �                      @        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    r@���Q��?             $@       �       �       	          ����?؇���X�?             @        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ���@@-�_ .�?�             g@       �       �                    @L@������?�            �f@       ������������������������       �        h             b@        �       �                   �s@؇���X�?            �A@       �       �                    c@XB���?             =@       ������������������������       �                     8@        �       �                   Pc@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?�q�q�?             @       �       �                   �d@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�b��	     h�h)h,K ��h.��R�(KK�KK��hb�B�
  �E$�~V�?�����?,������?u��QNG�?��9A��?'wc�#�?wwwwww�?""""""�?l�l��??�>��?              �?�$I�$I�?۶m۶m�?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?�������?�������?      �?                      �?              �?�$2���?���Id�?^Cy�5�?Q^Cy��?]t�E]�?F]t�E�?9��8���?�q�q�?      �?                      �?              �?B{	�%��?/�����?              �?      �?        �<�"h�?W'u_�?�������?�������?      �?        w�qG�?qG�wĽ?              �?�]�ڕ��?��+Q��?              �?ffffff�?�������?      �?        �������?�������?              �?�5��P�?(�����?              �?      �?        F]t�E�?/�袋.�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?TD�zaݵ?vW��SD�?�������?�������?{�G�z�?���Q��?              �?|���?>����?              �?�?�������?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?333333�?�������?�������?�������?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?��p�C�?n����{�?;�;��?O��N���?�1�K��?aw&��+�?      �?        UUUUUU�?UUUUUU�?              �?{�G�z�?���Q��?UUUUUU�?UUUUUU�?�A�A�?_�_��?�������?�������?              �?      �?      �?      �?                      �?              �?�؉�؉�?ى�؉��?              �?۶m۶m�?�$I�$I�?      �?                      �?              �?�������?�������?              �?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        S�n0�?�n0E>�?�5'���?�蕱���?�����?������?�������?KKKKKK�?�B!��?���{��?      �?      �?              �?F]t�E�?/�袋.�?      �?        �������?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?        ffffff�?333333�?      �?      �?      �?        KԮD�J�?jW�v%j�?      �?              �?      �?;�;��?b'vb'v�?l(�����?(������?      �?      �?      �?              �?      �?              �?      �?        F]t�E�?]t�E]�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?333333�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        S�n0E�?к����?�q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?GX�i���?�{a���?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�
HyhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK˅�h��B�2         �       
             �?
���P��?�           ��@              e                   �b@�n`���?            {@                                  �?,UP���?�             w@                                   b@     8�?"             P@                                  ]@X�<ݚ�?            �F@        ������������������������       �                     (@                                   �P@����e��?            �@@              	                    �?�q�q�?             >@        ������������������������       �                      @        
                           f@����X�?             <@                     	          `ff@z�G�z�?             9@                                 �^@�LQ�1	�?             7@                                   ]@���Q��?             @                                  @H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                  P`@�X�<ݺ?             2@       ������������������������       �                     *@                                   @M@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?�KM�]�?	             3@       ������������������������       �                     1@        ������������������������       �                      @               &                   �[@�˹�m��?�             s@                                   _@��<b���?             7@        ������������������������       �                     &@                !                    �?�q�q�?	             (@        ������������������������       �                      @        "       #                    �?�z�G��?             $@        ������������������������       �                     @        $       %       	             �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        '       *                   �Q@�@"�#�?�            �q@        (       )       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        +       `                    �Q@H�te�?�            `q@       ,       E                    �?�Xyd�B�?�            �p@        -       .                   `]@L紂P�?%            �I@        ������������������������       �                     1@        /       0                   @^@H�V�e��?             A@        ������������������������       �                      @        1       2                   �_@     ��?             @@        ������������������������       �                     @        3       8                    �L@���B���?             :@        4       5       	          ����?      �?             @        ������������������������       �                      @        6       7                    W@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        9       @                    �?ףp=
�?             4@       :       ?                   �l@�C��2(�?	             &@       ;       <       	             �?z�G�z�?             @        ������������������������       �                      @        =       >       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        A       D                   p`@�����H�?             "@        B       C                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        F       K                    �D@��6�.ӯ?�            @k@        G       H                    b@z�G�z�?             $@       ������������������������       �                     @        I       J                    �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        L       [       	          ����?���%�?�             j@        M       V                    �?�X�<ݺ?,             R@       N       O       	          433�? pƵHP�?              J@       ������������������������       �                     <@        P       Q                    @K@ �q�q�?             8@        ������������������������       �                     0@        R       U       	          ����?      �?              @        S       T                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        W       X                   �g@R���Q�?             4@        ������������������������       �                     (@        Y       Z                   �j@      �?              @        ������������������������       �                     @        ������������������������       �                     @        \       ]                    �?�|�l�?U             a@       ������������������������       �        8            �V@        ^       _                   �e@����?�?            �F@       ������������������������       �                     F@        ������������������������       �                     �?        a       b                   �[@�q�q�?             "@        ������������������������       �                     @        c       d                   `c@      �?             @       ������������������������       �                     @        ������������������������       �                     @        f       q                    �?      �?+            �P@        g       h                    m@      �?             <@        ������������������������       �                     &@        i       l       	          hff�?j���� �?
             1@        j       k                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        m       p                   �q@"pc�
�?             &@        n       o                    q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        r       �                    @�����?             C@       s       �                   @a@z�G�z�?             >@       t              	             @H%u��?             9@       u       z       	          ����?���}<S�?             7@        v       w       
             �?�q�q�?             @        ������������������������       �                     �?        x       y                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        {       ~                   �[@P���Q�?             4@        |       }       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             2@        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �       	          @33�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `f@      �?              @       �       �       	          @33�?      �?             @        ������������������������       �                     �?        �       �                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �f@R���Q�?�            �r@       �       �       	          ����?[�� ��?�            �r@       �       �                    �?�2<�Z��?�            �n@        �       �                   @Z@r�q��?-            �P@        ������������������������       �                      @        �       �                    �?     ��?,             P@        �       �                    �M@����X�?
             ,@       �       �                   �q@�C��2(�?             &@       ������������������������       �                     "@        �       �                   u@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �c@ףp=
�?"             I@       �       �                    �P@P�Lt�<�?             C@       ������������������������       �                    �B@        ������������������������       �                     �?        �       �                     H@�q�q�?	             (@       ������������������������       �                     @        �       �                   @`@z�G�z�?             @        ������������������������       �                     @        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�x�E~�?p            @f@        �       �                   0m@�C��2(�?             6@        �       �                   �a@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     2@        �       �                    @L@�(�Tw�?b            �c@       ������������������������       �        W             a@        �       �                    �L@�KM�]�?             3@        ������������������������       �                      @        ������������������������       �        
             1@        �       �                   pb@|��?���?%             K@       �       �                    �?r֛w���?             ?@        ������������������������       �                     @        �       �                    �?HP�s��?             9@       �       �                    �?z�G�z�?             $@        ������������������������       �                     @        �       �                   @^@����X�?             @        ������������������������       �                     �?        �       �                   �p@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �       �                    �?��<b���?             7@        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                    @M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    a@r�q��?             2@        �       �                     I@�z�G��?             $@        ������������������������       �                     @        �       �                    d@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  փmM���?>IY�8�?�c�1��?�9�s��?����7��?Y�B���?      �?     ��?r�q��?�q�q�?      �?        6�d�M6�?e�M6�d�?UUUUUU�?UUUUUU�?      �?        �$I�$I�?�m۶m��?�������?�������?Y�B��?��Moz��?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?��8��8�?              �?�������?�������?      �?                      �?      �?              �?              �?        (�����?�k(���?              �?      �?        ^Cy�5�?��P^Cy�?��Moz��?��,d!�?              �?�������?�������?      �?        333333�?ffffff�?              �?      �?      �?      �?                      �?�]�BO�?=Eԯ��?UUUUUU�?UUUUUU�?      �?                      �?���1O�?�_��?�f�P���?���U�?�������?�������?              �?ZZZZZZ�?iiiiii�?      �?              �?      �?              �?ى�؉��?��؉���?      �?      �?              �?      �?      �?              �?      �?        �������?�������?F]t�E�?]t�E�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?��p�?���A���?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ى�؉��?�;�;�?�q�q�?��8��8�?;�;��?'vb'vb�?              �?UUUUUU�?�������?              �?      �?      �?      �?      �?              �?      �?                      �?333333�?333333�?              �?      �?      �?      �?                      �?~?�������?              �?l�l��?��I��I�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?      �?      �?              �?ZZZZZZ�?�������?�������?UUUUUU�?      �?                      �?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?Q^Cy��?^Cy�5�?�������?�������?)\���(�?���Q��?ӛ���7�?d!Y�B�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?ffffff�?�������?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?�������?333333�?      �?              �?      �?      �?                      �?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?333333�?XY���a�?����Dx�?mާ�d�?.�u�y�?�������?UUUUUU�?              �?     ��?      �?�m۶m��?�$I�$I�?]t�E�?F]t�E�?      �?              �?      �?              �?      �?                      �?�������?�������?���k(�?(�����?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?      �?                      �?����G�?p�\��?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?        p��o���?�A�A�?      �?        �k(���?(�����?              �?      �?        	�%����?{	�%���?�B!��?���{��?      �?        {�G�z�?q=
ףp�?�������?�������?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?                      �?��,d!�?��Moz��?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���]hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK˅�h��B�2         v                    �?R������?�           ��@              A       
             �?&���7��?           �{@                      	          ����?>��"��?n            �e@                                   �?�[|x��?             �O@                                  �?4?,R��?             B@        ������������������������       �        	             3@                                  @b@�t����?	             1@        ������������������������       �                     $@        	                           �?����X�?             @        
                           �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@               :                   Xr@      �?N            �[@                                 �\@��V�I��?B            �W@        ������������������������       �                     ,@                                   �?�Q����?7             T@                                   �K@�θ�?             :@                                  @I@�}�+r��?             3@                                  �G@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@                                  m@����X�?             @        ������������������������       �                      @        ������������������������       �                     @               7                     P@�5��?(             K@              "       
             �?�G��l��?              E@                                  �j@�����H�?             "@        ������������������������       �                     @                !                    d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        #       *                   �l@���|���?            �@@       $       )                    �N@     ��?             0@       %       &                    W@���|���?             &@        ������������������������       �                     @        '       (                   �a@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        +       2                    �K@@�0�!��?             1@        ,       -                   �n@���Q��?             @        ������������������������       �                      @        .       /                   �c@�q�q�?             @        ������������������������       �                     �?        0       1                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       6       	          ����?�8��8��?             (@        4       5                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        8       9                   �c@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ;       @                    �?     ��?             0@       <       ?                    b@�z�G��?             $@       =       >       	          pff@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        B       O                    c@�NJa&��?�            �p@        C       N                    �?r�q��?             8@       D       E                    �?     ��?	             0@        ������������������������       �                     �?        F       G                   `Y@�r����?             .@        ������������������������       �                     �?        H       I                    �?@4և���?             ,@        ������������������������       �                     "@        J       K                    @G@z�G�z�?             @        ������������������������       �                      @        L       M                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        P       Q                   @i@ @|���?�            �n@        ������������������������       �        (            �P@        R       s                    c@������?l            @f@       S       T                   pi@�q�Y��?g            @e@        ������������������������       �                     �?        U       p                    @ 
��р�?f             e@       V       ]                    �I@�6,r➷?d            �d@       W       X                    �?��F�D�?8            �X@        ������������������������       �                     C@        Y       \                    �?�]0��<�?"            �N@        Z       [                   `\@؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                    �G@        ^       c                    @J@�C��2(�?,            �P@        _       b                    �?z�G�z�?
             .@        `       a                   �l@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        d       o                   �c@�IєX�?"            �I@       e       f                     L@     ��?             @@        ������������������������       �                     (@        g       h                   Hp@R���Q�?             4@        ������������������������       �                      @        i       j                    �L@      �?             (@        ������������������������       �                      @        k       l                   ps@ףp=
�?             $@       ������������������������       �                     @        m       n                   �v@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        q       r                   Pl@      �?             @        ������������������������       �                      @        ������������������������       �                      @        t       u                   �c@      �?              @       ������������������������       �                     @        ������������������������       �                     @        w       �       
             �?�6hܟo�?�            Pr@       x       �                    �?�}#���?�             o@        y       |       	          ����?¦	^_�?             ?@        z       {                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        }       �                   �k@�J�4�?             9@        ~                           a@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �q@ףp=
�?             4@        ������������������������       �                     "@        �       �                   @_@"pc�
�?             &@        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       �       �                   �r@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��Ujѡ�?�            @k@       �       �                    �M@P4�!*ͯ?y            `g@       �       �                    �?Hn�.P��?Q             _@       �       �                   �i@���.�6�?=             W@        ������������������������       �                     =@        �       �                   �Z@�����?,            �O@        ������������������������       �                     �?        �       �                   �\@6uH���?+             O@        �       �                   `[@�<ݚ�?             2@       �       �                   �W@@4և���?
             ,@        ������������������������       �                     @        �       �                    �?؇���X�?             @       ������������������������       �                     @        �       �                   (q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �k@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   0c@`���i��?             F@       ������������������������       �                     E@        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @@        ������������������������       �        (            �O@        �       �                   0b@�n`���?             ?@       �       �                    �?H%u��?             9@        ������������������������       �                      @        �       �                   @^@�nkK�?             7@        �       �                   �\@      �?              @        ������������������������       �                     @        �       �                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        �       �                   c@      �?             @        ������������������������       �                      @        �       �                   ``@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �\@d�
��?              F@        ������������������������       �                     @        �       �                   �j@��
ц��?            �C@        �       �                    �?�θ�?             *@       �       �                   �`@      �?
             (@        �       �                    �O@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    n@�	j*D�?             :@        ������������������������       �                      @        �       �                    �?X�<ݚ�?             2@        ������������������������       �                     @        �       �                     R@�q�q�?	             (@       �       �                     K@���Q��?             $@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @`@���Q��?             @        ������������������������       �                      @        �       �       	          `ff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��*��?5��j���?͎Z���?e�J��?��R�O2�?�����?EQEQ�?]�u]�u�?r�q��?�8��8��?              �?�������?�������?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?r1����?G}g����?              �?�������?ffffff�?ى�؉��?�؉�؉�?�5��P�?(�����?�q�q�?�q�q�?      �?                      �?      �?        �$I�$I�?�m۶m��?      �?                      �?/�����?h/�����?��y��y�?1�0��?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?]t�E]�?      �?      �?F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?              �?      �?              �?        �������?ZZZZZZ�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?UUUUUU�?�������?              �?      �?              �?      �?ffffff�?333333�?      �?      �?      �?                      �?              �?      �?        ~5&��?IT�n�?UUUUUU�?UUUUUU�?      �?      �?              �?�������?�?              �?n۶m۶�?�$I�$I�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?"XG��)�?�}�K�`�?      �?        ؽ�u�{�?B�P�"�?�������?�������?              �?	j*D�?�n_Y�K�?s�,��r�?�0�Ө?j�J�Z�?[�R�֯�?      �?        \2�h��?;ڼOqɠ?۶m۶m�?�$I�$I�?              �?      �?              �?        ]t�E�?F]t�E�?�������?�������?�������?333333�?              �?      �?              �?        �?�?      �?      �?      �?        333333�?333333�?      �?              �?      �?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?              �?      �?      �?                      �?�L��Y�?���Z�i�?4u~�!��?Y1P�M�?�RJ)���?��Zk���?�������?UUUUUU�?      �?                      �?{�G�z�?�z�G��?�������?333333�?              �?      �?        �������?�������?              �?F]t�E�?/�袋.�?      �?        �������?�������?�$I�$I�?۶m۶m�?      �?                      �?              �?��A��.�?��p=�?n�ʄm�?�>V�'��?�c�1ƨ?t�9�s�?Y�B��?���7���?              �?�a�a�?=��<���?      �?        ��RJ)��?k���Zk�?�q�q�?9��8���?�$I�$I�?n۶m۶�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?      �?              �?      �?        F]t�E�?F]t�E�?              �?      �?      �?      �?                      �?              �?              �?�c�1��?�9�s��?���Q��?)\���(�?      �?        d!Y�B�?�Mozӛ�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?              �?      �?              �?      �?        �.�袋�?�袋.��?              �?�;�;�?�؉�؉�?�؉�؉�?ى�؉��?      �?      �?      �?      �?      �?                      �?              �?              �?vb'vb'�?;�;��?      �?        r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?�������?333333�?�������?�������?      �?                      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�;hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKم�h��B@6         �                    �?�r,��?�           ��@              Y       	             �?Ή�Bk��?           �z@                                 �\@�θ�?�            �u@                      
             �?Z�K�D��?            �G@                                  �?      �?             @@                                   @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        	              	          033�?$�q-�?             :@       
                           �?�nkK�?             7@                                 @^@��S�ۿ?
             .@                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @                                  �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�r����?	             .@       ������������������������       �                     (@                                  �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �c@���a��?�             s@                      
             �?J�8���?             =@        ������������������������       �                     @                      
             �?�+e�X�?             9@       ������������������������       �        	             1@                      	             �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        !       @       
             �?䦳	�R�?�            0q@        "       ?                    @N@�G\�c�?'            @P@       #       >                   @a@��o	��?"             M@       $       7                   p@�E��
��?             J@       %       ,       	          ����?����X�?            �A@        &       +                    �?      �?             ,@       '       (                    �?�z�G��?             $@        ������������������������       �                      @        )       *                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        -       .                   l@؇���X�?             5@        ������������������������       �                     $@        /       0                    �?���!pc�?             &@        ������������������������       �                     @        1       2                    �F@      �?             @        ������������������������       �                      @        3       4       
             �?      �?             @        ������������������������       �                      @        5       6                    @J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        8       ;                   `r@ҳ�wY;�?	             1@       9       :                    `@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        <       =       	             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        A       H                    �L@�Ń��̧?�            @j@       B       G                    �?@�����?p             e@        C       F                   0k@P�Lt�<�?             C@        D       E       	          ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �        Y            ``@        I       R                    �?������?            �D@        J       K                   �b@z�G�z�?	             .@        ������������������������       �                      @        L       Q       	          ����?և���X�?             @       M       N                   @d@�q�q�?             @        ������������������������       �                     �?        O       P                   �r@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        S       X                   �`@ ��WV�?             :@        T       U                    �?      �?              @        ������������������������       �                     �?        V       W                    @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             2@        Z       {       
             �?���!pc�?4            @S@       [       n                   �b@���*�?(             N@       \       c                    �?X�EQ]N�?            �E@        ]       b                    �?      �?              @       ^       a                    �?r�q��?             @       _       `                   �_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        d       e       	          ����? >�֕�?            �A@        ������������������������       �                     2@        f       i                   �]@�t����?             1@        g       h                   �[@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        j       k                    �?@4և���?	             ,@        ������������������������       �                      @        l       m                   pl@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        o       z                   `d@ҳ�wY;�?             1@       p       u                   �^@��
ц��?	             *@        q       t                   �c@؇���X�?             @        r       s                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        v       y                   �c@r�q��?             @        w       x                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        |       }                    �?j���� �?             1@       ������������������������       �                     "@        ~       �                    �M@      �?              @               �                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?0�����?�             s@       �       �                    @G@أ����?�            �n@        �       �                    �?���!pc�?            �@@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?PN��T'�?             ;@       �       �                    b@�����?             5@       ������������������������       �                     2@        �       �                    _@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	             �?�q�q�?             @        ������������������������       �                      @        �       �                   �l@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �d@� Λ��?�            �j@       �       �       
             �?HH�^'д?�            �j@       �       �                   @^@�w��3(�?t            �g@        �       �                    �I@      �?             8@        �       �                   �\@�q�q�?             @        ������������������������       �                     @        �       �                    Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?�X�<ݺ?             2@        �       �                    �K@r�q��?             @        ������������������������       �                     @        �       �                   @[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   `\@�Sa��?f            �d@        �       �                     R@�.ߴ#�?&            �N@       �       �                    `@(;L]n�?%             N@        �       �       	          ����?؇���X�?             @       �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?�O4R���?"            �J@        �       �                   @a@r�q��?             @        ������������������������       �                      @        �       �                    �?      �?             @       �       �                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �G@        ������������������������       �                     �?        ������������������������       �        @            �Z@        �       �       	             �?؇���X�?             5@        �       �                   �^@      �?             @        ������������������������       �                      @        �       �                     N@      �?             @        �       �                   �h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                      @        �       �       
             �? 1_#�?#            �M@       �       �                   �i@     ��?             H@        ������������������������       �                     2@        �       �                   �\@�z�G��?             >@        ������������������������       �                     @        �       �                   Pk@���B���?             :@        �       �                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �s@�C��2(�?             6@       �       �                   `b@P���Q�?             4@       ������������������������       �                     ,@        �       �                     P@r�q��?             @        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?"pc�
�?             &@       ������������������������       �                     @        �       �                    �K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �292ȯ�?�f����?
�N]���?�bEi|�?ى�؉��?�؉�؉�?]AL� &�?R�٨�l�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?�؉�؉�?d!Y�B�?�Mozӛ�?�?�������?�������?�������?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�k(���?��P^Cy�?|a���?�rO#,��?      �?        ���Q��?R���Q�?              �?      �?      �?      �?                      �?G�kĿF�?���ʽ?S+�R+��?[��Z���?���{�?������?;�;��?��؉���?�m۶m��?�$I�$I�?      �?      �?ffffff�?333333�?              �?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?        F]t�E�?t�E]t�?      �?              �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?�������?�������?UUUUUU�?�������?              �?      �?        �������?�������?              �?      �?                      �?      �?        ��<��<�?�a�a�?��
ц��?ݾ�z�<x?���k(�?(�����?      �?      �?      �?                      �?      �?              �?        �|����?������?�������?�������?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?              �?O��N���?;�;��?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?        t�E]t�?F]t�E�?wwwwww�?""""""�?qG�wĽ?w�qG�?      �?      �?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        �A�A�?��+��+�?              �?�?<<<<<<�?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�؉�؉�?�;�;�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?�������?ZZZZZZ�?      �?              �?      �?      �?      �?              �?      �?                      �? u�uʿ?\�\��?�KA���?���h�?t�E]t�?F]t�E�?�������?UUUUUU�?      �?                      �?h/�����?&���^B�?�a�a�?=��<���?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        7��XQ�?�L�w�Z�?�琚`��?��V�9��?kP<�q�?�:,���?      �?      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?��8��8�?UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?7Āt,e�?��[��l�?XG��).�?�K�`m�?�?�������?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?�x+�R�?:�&oe�?UUUUUU�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?      �?              �?      �?              �?                      �?      �?        ��c+���?	N�<�?      �?      �?              �?333333�?ffffff�?      �?        ى�؉��?��؉���?      �?      �?      �?                      �?F]t�E�?]t�E�?�������?ffffff�?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?/�袋.�?F]t�E�?      �?              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ� �thG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@,         b                    �?�[��N�?�           ��@                                  P@f�B���?           �y@                                   @N@`����x�?I            �\@                                  �?`-�I�w�?0             S@                      
             �?r�q��?             >@       ������������������������       �                     2@                                  @b@�q�q�?	             (@                     	          @33�?�z�G��?             $@        	       
                    @I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                      	             �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     G@        ������������������������       �                     C@               5       	          pff�?0,Tg��?�            `r@               "       
             �?���o� �??            �Y@                                  pb@�z�G��?             D@                                  \@r�q��?             >@                                   �?X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @                      	          ����?���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?               !                   �d@�z�G��?             $@                                   �?      �?              @                     	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        #       $                   �b@���N8�?'            �O@       ������������������������       �                     ?@        %       .                    �?     ��?             @@       &       -       	          ����?�t����?             1@       '       *                    �L@؇���X�?             ,@       (       )                   �c@�8��8��?
             (@        ������������������������       �                     �?        ������������������������       �        	             &@        +       ,                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        /       0                    �?�q�q�?             .@        ������������������������       �                     @        1       2                    p@r�q��?             (@        ������������������������       �                     @        3       4                   `e@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        6       M       	          ����?(�_���?{            �g@        7       8       
             �?�iʫ{�?!            �J@        ������������������������       �                      @        9       @                    �?L紂P�?             �I@        :       ;                   �^@      �?              @        ������������������������       �                     �?        <       =                     L@����X�?             @        ������������������������       �                     @        >       ?                   �q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        A       L                   �e@�ʈD��?            �E@       B       C                   ``@@4և���?             E@       ������������������������       �                     <@        D       G                   �`@d}h���?             ,@        E       F                     J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        H       I       
             �?�C��2(�?             &@       ������������������������       �                      @        J       K                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        N       a                   �d@p��%���?Z            @a@       O       ^                    `R@ 7���B�?X            �`@       P       Q                   �Z@�z�N��?U            ``@        ������������������������       �                     �?        R       S                   `_@ ����?T            @`@       ������������������������       �        1             R@        T       W                   `i@XB���?#             M@        U       V                   �\@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        X       Y                    @P@�O4R���?            �J@       ������������������������       �                    �H@        Z       ]       	          ���@      �?             @       [       \                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        _       `                   �p@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        c       �                    �?*��In�?�            `t@       d       �                    @L@�A����?�            �p@       e       �                    @P���+�?�            �h@       f       �       
             �?(�_���?}            �g@        g       l                    �G@`��}3��?             �J@        h       k                    @B@�����?             5@        i       j       	              @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             1@        m       �                   ``@     ��?             @@       n       u       
             �?�z�G��?             4@        o       p                    �?ףp=
�?             $@        ������������������������       �                     @        q       t                   Pm@؇���X�?             @       r       s                    ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        v       w                   `]@      �?             $@        ������������������������       �                     @        x       y                    �?����X�?             @        ������������������������       �                     @        z                          �^@      �?             @       {       |       	          ����?�q�q�?             @        ������������������������       �                     �?        }       ~       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             (@        ������������������������       �                      @        �       �                   �d@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �        ]            @a@        �       �       	          ����?      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?�\����?)            �P@       �       �                   �c@�<ݚ�?             B@       �       �                   `V@�c�Α�?             =@        ������������������������       �                     @        �       �                    c@���B���?             :@       �       �                    X@      �?             8@        ������������������������       �                     �?        �       �                   �s@���}<S�?             7@       �       �                    �?���7�?             6@       ������������������������       �                     4@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?�������?             >@        ������������������������       �                      @        �       �                   @b@�>4և��?             <@       �       �                    �?HP�s��?             9@       �       �                     Q@ �q�q�?             8@       ������������������������       �        
             4@        �       �                   �n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����5�?"            �N@        ������������������������       �                      @        �       �                   �_@�T`�[k�?            �J@       ������������������������       �                     >@        �       �                   �f@
;&����?             7@       �       �                   �n@p�ݯ��?             3@       �       �                   `Z@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        �       �                   0`@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  B~�9�J�?�@c�Z�?�������?�������?Lg1��t�?��,����?y�5�װ?Q^Cy��?UUUUUU�?�������?              �?�������?�������?333333�?ffffff�?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?                      �?              �?1�0��?�y��y��?r^�	��?C���?333333�?ffffff�?UUUUUU�?�������?�q�q�?r�q��?              �?      �?        �a�a�?��y��y�?              �?      �?        ffffff�?333333�?      �?      �?      �?      �?              �?      �?              �?                      �?�a�a�?��y��y�?      �?              �?      �?�������?�������?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?              �?�������?333333�?              �?      �?        �qɶ?�Q�}�&�?�琚`��?
�[���?      �?        �������?�������?      �?      �?      �?        �$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        �}A_з?A_���?�$I�$I�?n۶m۶�?              �?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        ہ�v`��?�g��%�?h/�����?	�%����?ձ�6Ls�?qBJ�eD�?      �?         �����? �����?              �?�{a���?GX�i���?�������?�������?      �?                      �?�x+�R�?:�&oe�?              �?      �?      �?      �?      �?      �?                      �?              �?      �?      �?              �?      �?              �?        |��¬�?�ɀz��?T�ѯz�?үz�@�?���/M�?�Q7���?�Q�}�&�?�qɶ?�琚`��?M0��>��?=��<���?�a�a�?      �?      �?      �?                      �?      �?              �?      �?ffffff�?333333�?�������?�������?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?�m۶m��?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?      �?      �?        �������?�������?              �?      �?              �?              �?      �?              �?      �?        ���>��?>����?9��8���?�q�q�?5�rO#,�?�{a���?              �?��؉���?ى�؉��?      �?      �?              �?ӛ���7�?d!Y�B�?�.�袋�?F]t�E�?      �?              �?      �?              �?      �?                      �?              �?      �?        �������?�������?      �?        �m۶m��?�$I�$I�?{�G�z�?q=
ףp�?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?              �?        ������?��).��?      �?        "5�x+��?���!5��?              �?Y�B��?�Mozӛ�?^Cy�5�?Cy�5��?;�;��?;�;��?              �?      �?        UUUUUU�?�������?      �?                      �?              �?�t�bub�      hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��1hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKÅ�h��B�0         x       
             �?"�\�&U�?�           ��@              K                    �?�^о�?           p{@                                   �?�H�a��?l            @e@                     	            �?��{H�?<            �U@        ������������������������       �                     =@                                  �a@>���Rp�?(             M@                     	          ����?p�ݯ��?             C@               	                    �?������?             1@        ������������������������       �                     @        
                          pd@�q�q�?
             (@                                 P`@      �?              @                                  `@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                  �]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   @O@���N8�?             5@       ������������������������       �        	             0@                                   �?z�G�z�?             @        ������������������������       �                     @                                  @\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@               F                    �?��q7L��?0            �T@              #                   �h@(ǯt��?+            �R@               "                    �Q@�θ�?             *@                                 �f@�C��2(�?             &@        ������������������������       �                     @                !                   @`@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        $       C                    �?Nd^����?$            �N@       %       &                   `X@r�z-��?             �J@        ������������������������       �                      @        '       *       
             �?�\�u��?            �I@        (       )                    �I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        +       2                    �?(���@��?            �G@        ,       -                   0q@ףp=
�?             4@       ������������������������       �        
             .@        .       1                    @L@���Q��?             @       /       0                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        3       4                   `]@|��?���?             ;@        ������������������������       �                      @        5       >                    �?� �	��?             9@        6       9                    _@      �?             (@        7       8       	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        :       ;                    d@����X�?             @        ������������������������       �                      @        <       =                   p@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ?       B       	          ���@�n_Y�K�?             *@       @       A                   0a@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        D       E                    r@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        G       J                    @K@�����H�?             "@        H       I                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        L       W                    �?|�db���?�            �p@        M       P                    @G@�k�'7��?!            �L@        N       O                   0b@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        Q       V                    @`�q�0ܴ?            �G@       R       U                   �\@��<b�ƥ?             G@        S       T                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     F@        ������������������������       �                     �?        X       w                    �?HH�^'д?�            �j@       Y       t                   �b@p��D׀�?a            �c@       Z       ]                   @Z@P-�T6��?]            �b@        [       \                   Pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ^       q                   �u@hڛ�ʚ�?[            �b@       _       p       	          ����?@��8��?W             b@       `       o                    �? 7���B�?0            @T@       a       b                   Pe@���N8�?&            �O@        ������������������������       �                     6@        c       h                   �Z@��p\�?            �D@        d       g                    @N@؇���X�?             ,@       e       f                   0j@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        i       j                    _@ 7���B�?             ;@        ������������������������       �                     (@        k       l       	          ����?��S�ۿ?             .@       ������������������������       �                     &@        m       n                   Ph@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             2@        ������������������������       �        '            �O@        r       s       	          ����?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        u       v                     D@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        "             K@        y       �                   @E@Vi1�;$�?�            pr@        z       �       	          ����?д>��C�?             =@        {       |                    �?���Q��?             @        ������������������������       �                      @        }       ~                   �a@�q�q�?             @        ������������������������       �                     �?               �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@�8��8��?             8@       ������������������������       �        	             *@        �       �                   a@"pc�
�?             &@        ������������������������       �                     �?        �       �       	          hff�?ףp=
�?             $@        �       �                    c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?`�t欝�?�            �p@        �       �                    �?��It��?1            �S@        �       �                    �?�f7�z�?             =@       �       �                    �?      �?             0@       �       �                    �?�q�q�?             "@        ������������������������       �                     �?        �       �                    @J@      �?              @       �       �                   �o@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @K@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �I@ףp=
�?#             I@       ������������������������       �                     =@        �       �                   pc@���N8�?             5@       �       �       	          433�?@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        �       �                   �]@և���X�?             @        ������������������������       �                     @        �       �                   �i@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    c@��R�x��?w            `g@       �       �                   �^@XB���?n            �e@       �       �                    �? }�Я��?8            @V@       ������������������������       �        !             L@        �       �                    @H@Pa�	�?            �@@       ������������������������       �                     2@        �       �                     I@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                   Pd@�IєX�?6            @U@       �       �                   �s@��ϭ�*�?$             M@       �       �                    _@ �h�7W�?             �J@        ������������������������       �                      @        �       �                   �c@���J��?            �I@       ������������������������       �                     H@        �       �                   pn@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���Q��?             @        �       �                   Hv@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                    �?8�Z$���?	             *@        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  ��j��`�?:�J;�O�?*���H�?�}�ƭ�?TTTTTT�?�������?/�I���?���C���?              �?GX�i���?�i��F�?Cy�5��?^Cy�5�?xxxxxx�?�?      �?        UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?�a�a�?��y��y�?              �?�������?�������?              �?      �?      �?              �?      �?                      �?��FS���?��\V��?���g��?S�n0E�?�؉�؉�?ى�؉��?F]t�E�?]t�E�?              �?UUUUUU�?�������?      �?                      �?      �?        �u�y���?���:�?����!�?�琚`��?              �?�������?�?      �?      �?              �?      �?        W�+���?R�٨�l�?�������?�������?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        {	�%���?	�%����?              �?�Q����?)\���(�?      �?      �?�������?�������?      �?                      �?�$I�$I�?�m۶m��?              �?�������?333333�?      �?                      �?;�;��?ى�؉��?�q�q�?�q�q�?      �?                      �?              �?      �?      �?              �?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?�Q���?�ĵb��?Lg1��t�?-����b�?�������?�������?              �?      �?        W�+�ɥ?��F}g��?d!Y�B�?��7��M�?      �?      �?              �?      �?                      �?      �?        �琚`��?��V�9��?T:�g *�?[܄�]-�?�`Q�(X�?���t}��?      �?      �?      �?                      �?7`��c.�?�y����?UUUUUU�?UUUUUU�?h/�����?	�%����?�a�a�?��y��y�?              �?��+Q��?�]�ڕ��?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?      �?                      �?      �?        h/�����?	�%����?              �?�?�������?              �?      �?      �?      �?                      �?              �?              �?�������?333333�?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?                      �?�B��r$�?����5n�?|a���?a���{�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?F]t�E�?/�袋.�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?A�d�?���7G߼?-n����?�#{���?a���{�?O#,�4��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?�������?              �?      �?              �?              �?        ;�;��?;�;��?      �?                      �?�������?�������?      �?        �a�a�?��y��y�?n۶m۶�?�$I�$I�?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?      �?              �?      �?        ��rD���?�и[�?GX�i���?�{a���?�я~���?p�\��?      �?        |���?|���?      �?        �������?�?              �?      �?        �?�?����=�?|a���?��sHM0�?"5�x+��?              �?______�?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�JIhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@(         j       
             �?�_y���?�           ��@                                 0b@D>�Q�?            z@                                  @^@ȑ����?G            @]@                                  �?$Q�q�?'            �O@                                   �?8�Z$���?             :@       ������������������������       �                     3@                      	          `ff�?և���X�?             @              	                   �T@���Q��?             @        ������������������������       �                      @        
                           @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �B@        ������������������������       �                      K@               E                    �?�><Ym}�?�            �r@                                 �Z@4��?�?�             j@                      	          ����?�q�q�?             @        ������������������������       �                     �?                                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               2       	          ����?���(��?�            �i@                                   �?�M���?-             Q@                                   �M@�eP*L��?
             &@        ������������������������       �                     @        ������������������������       �                     @               %                    �?�S����?#            �L@               $                    �?�eP*L��?
             &@                                  �J@���Q��?	             $@       ������������������������       �                     @                #                   �_@z�G�z�?             @        !       "                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        &       '                    @K@���}<S�?             G@       ������������������������       �                     5@        (       /       	          ����?�J�4�?             9@       )       .                    �?�C��2(�?
             6@       *       +       	          ����?r�q��?             (@        ������������������������       �                     @        ,       -                   �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        0       1                    Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        3       4                   �c@`Y����?T             a@        ������������������������       �                     �?        5       <                    \@ ��ʻ��?S             a@        6       7                   `_@r�q��?             @        ������������������������       �                      @        8       ;                   �`@      �?             @        9       :                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        =       D                    _@��G^�C�?N            @`@        >       C                    �J@�IєX�?	             1@       ?       B                   �p@      �?              @       @       A                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �        E            @\@        F       G                    @G@rѱ�D��?:            �V@        ������������������������       �                     "@        H       M                    �?�W����?2            �T@        I       J                   `X@�KM�]�?             3@        ������������������������       �                     �?        K       L                   `c@�X�<ݺ?
             2@       ������������������������       �        	             1@        ������������������������       �                     �?        N       Y                   a@b����?'            �O@        O       R                    �?HP�s��?             9@        P       Q                    `P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       T                   �]@�nkK�?             7@       ������������������������       �                     (@        U       V                    �?�C��2(�?             &@       ������������������������       �                     @        W       X                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       ]                    @I@�\��N��?             C@        [       \                   0f@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ^       i                   Xq@l��
I��?             ;@       _       h                    `P@�q�q�?             8@       `       g                    �N@�㙢�c�?             7@       a       f       	             @������?
             1@       b       c                   0o@@4և���?             ,@       ������������������������       �                     (@        d       e       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        k       �       	             �?���U�?�            �s@       l       �                    �?��L��?�            �q@        m       x                   @E@����"�?8            �U@        n       q                    �M@�E��ӭ�?             2@       o       p                   `[@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        r       s                   Pa@�q�q�?             @        ������������������������       �                     �?        t       w       	             �?z�G�z�?             @       u       v                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        y       �                    �?(���X�?,            @Q@       z       {                   �b@r�����?!            �J@       ������������������������       �                     =@        |       �                    @J@�q�q�?             8@        }       �                   �_@�q�q�?             (@       ~                           �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    s@r�q��?             (@       �       �                    \@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �?      �?             0@        ������������������������       �                     @        �       �                   �b@�θ�?	             *@       �       �                    n@���Q��?             @        ������������������������       �                      @        �       �                    @J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �_@�a�O�?y            @h@        �       �       	          ����?XB���?             =@       ������������������������       �                     <@        ������������������������       �                     �?        �       �                   �i@��ϩ}��?e            �d@        �       �                    �L@�O4R���?!            �J@       ������������������������       �                     I@        �       �                   @b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        D             \@        �       �                    �?���"͏�?            �B@        �       �                   `T@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   pb@�r����?             >@       ������������������������       �                     :@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B
  V�.�#��?աh6n��?vb'vb'�?b'vb'v�?���?��~���?AA�?~��}���?;�;��?;�;��?              �?�$I�$I�?۶m۶m�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?���A�?�H����?ى�؉��?�N��N��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        z�gaz�?1=ӳ0�?<<<<<<�?�������?t�E]t�?]t�E�?      �?                      �?^Cy�5�?(������?]t�E�?t�E]t�?�������?333333�?              �?�������?�������?      �?      �?              �?      �?              �?              �?        d!Y�B�?ӛ���7�?              �?{�G�z�?�z�G��?F]t�E�?]t�E�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�d�*al�?�,���L�?      �?        �?�������?UUUUUU�?�������?              �?      �?      �?      �?      �?              �?      �?                      �? ����?�����?�?�?      �?      �?      �?      �?              �?      �?                      �?              �?              �?���?��=��=�?      �?        p>�cp�?��|���?�k(���?(�����?              �?��8��8�?�q�q�?      �?                      �?�eY�eY�?5M�4M��?{�G�z�?q=
ףp�?      �?      �?              �?      �?        d!Y�B�?�Mozӛ�?              �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?y�5���?�5��P�?F]t�E�?]t�E�?              �?      �?        Lh/����?h/�����?UUUUUU�?�������?�7��Mo�?d!Y�B�?xxxxxx�?�?n۶m۶�?�$I�$I�?      �?              �?      �?      �?                      �?              �?      �?                      �?              �?a��}��?~�	�[�?����?�\���?	�=����?�i��F�?r�q��?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?              �?      �?              �?        l�ځ��?)�3J���?Dj��V��?�V�9�&�?      �?        �������?�������?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?                      �?      �?        �������?UUUUUU�?]t�E�?F]t�E�?              �?      �?                      �?      �?      �?      �?        �؉�؉�?ى�؉��?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �? tT����?����?GX�i���?�{a���?      �?                      �?Ο��Y��?�0��x?:�&oe�?�x+�R�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        *�Y7�"�?v�)�Y7�?�m۶m��?�$I�$I�?              �?      �?        �?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��NhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�=         �                    �?�+	G�?�           ��@                                 �_@��j�+i�?           �z@                                   �N@�����?-             Q@                                 @E@�����?             E@                                 �a@$�q-�?            �C@                     
             �?R���Q�?             4@       ������������������������       �                     *@                                  @_@և���X�?             @       	                            I@z�G�z�?             @        
                           ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@                      
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �?$��m��?             :@                                   �?      �?              @                                  @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?�����H�?
             2@       ������������������������       �                     .@                                  �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               g                    @L@����s�?�            @v@              <                    �?6C�d�?�            �o@                ;                    �?     ��?+             P@       !       (       
             �?X�Cc�?%             L@        "       '                    �F@������?             1@        #       $                    �?z�G�z�?             @        ������������������������       �                     @        %       &       	          @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        )       *                    �?:�&���?            �C@        ������������������������       �                      @        +       4                   �l@��a�n`�?             ?@        ,       /                    �?X�Cc�?
             ,@        -       .                    @F@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        0       3                   �_@���Q��?             $@        1       2                   �b@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        5       :                   @_@�t����?
             1@        6       7                   �[@����X�?             @        ������������������������       �                     @        8       9                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        =       `       	          033�?��8��)�?v            �g@       >       ?                   pa@�����?r            �f@        ������������������������       �                     ?@        @       G                    �G@ghډC�?]            �b@       A       B                    �?`��F:u�?7            �U@        ������������������������       �                     ;@        C       D                   �a@��S�ۿ?#             N@        ������������������������       �                      @        E       F                   �c@XB���?"             M@        ������������������������       �                      @        ������������������������       �        !             L@        H       K                    g@؇���X�?&            �O@        I       J                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        L       W                    @I@�^����?$            �M@        M       V       	          ����?      �?             (@       N       S                    �?      �?              @       O       P                   �e@r�q��?             @        ������������������������       �                     @        Q       R                   0f@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        T       U                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        X       _       
             �?`Ql�R�?            �G@        Y       ^                   @c@�8��8��?             (@        Z       [                   �b@z�G�z�?             @        ������������������������       �                      @        \       ]       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �A@        a       b                    �?����X�?             @        ������������������������       �                     �?        c       f       	             @r�q��?             @       d       e                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        h       �       
             �?��
ц��?G             Z@       i       v                    �?J��D��?$             K@       j       u                   �d@�+$�jP�?             ;@       k       n                   p`@H%u��?             9@        l       m                   �\@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        o       t       	          ����?�}�+r��?             3@        p       s                    �?      �?              @        q       r                    �M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                      @        w       x       	          ����?X�<ݚ�?             ;@        ������������������������       �                     "@        y       �                    �?�q�q�?             2@       z       {                   �Z@؇���X�?
             ,@        ������������������������       �                     �?        |                          �`@$�q-�?	             *@       }       ~                   �`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �b@H.�!���?#             I@       �       �                    @ףp=
�?             >@       �       �                   Hp@�nkK�?             7@       ������������������������       �        
             0@        �       �                   pp@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                   Pp@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �g@���Q��?             4@        ������������������������       �                     @        �       �                    �?      �?             0@       �       �                    �N@�<ݚ�?             "@       �       �                   �e@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �i@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �Y@�jqL���?�            `s@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@ a�ox��?�            s@       �       �                    @R@�8��8��?�            @q@       �       �                    �?t�e�í�?�            �p@       �       �                    f@�P�U`��?z            `h@       �       �                   �s@��y� �?s            @g@       �       �       
             �?p��@���?g            @e@       �       �                    `@��F��?_            `c@        �       �                    �O@�t����?            �I@       �       �                    �?���}<S�?             G@       �       �                    �K@�7��?            �C@       ������������������������       �                     7@        �       �                    �?      �?	             0@       �       �                   �\@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @]@����X�?             @        �       �                    @K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   p`@���Q��?             @        ������������������������       �                      @        �       �                   �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �K@ pƵHP�?C             Z@        �       �                    �?���N8�?             E@        �       �       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @K@P�Lt�<�?             C@       ������������������������       �                     ?@        �       �                   �[@؇���X�?             @        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        '             O@        �       �       	          ����?������?             .@        ������������������������       �                     @        ������������������������       �                     &@        �       �                   ``@      �?             0@        �       �                    Z@X�<ݚ�?             "@        ������������������������       �                      @        �       �                   �\@և���X�?             @        ������������������������       �                      @        �       �                     M@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                   �a@      �?             @        ������������������������       �                      @        �       �                    �?      �?             @       �       �                     L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   a@ �й���?,            @R@       ������������������������       �        #             M@        �       �                   @m@��S�ۿ?	             .@       ������������������������       �                     $@        �       �                   c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �n@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                   0m@П[;U��?             =@        �       �                     G@ףp=
�?             $@        �       �                     D@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���y4F�?             3@       �       �                    @E@������?	             .@        ������������������������       �                     �?        �       �                    e@d}h���?             ,@       �       �                    @N@ףp=
�?             $@       ������������������������       �                     @        �       �                    �O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   pf@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  ��C�l�?z?+^���?~�	�[�?��sH�?xxxxxx�?�������?�a�a�?=��<���?;�;��?�؉�؉�?333333�?333333�?              �?۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        vb'vb'�?�N��N��?      �?      �?      �?      �?      �?                      �?      �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?�"�E�?�u�{���?˲,˲,�?�4M�4M�?      �?      �?%I�$I��?�m۶m��?�?xxxxxx�?�������?�������?      �?              �?      �?              �?      �?                      �?�A�A�?�o��o��?      �?        �c�1��?�s�9��?%I�$I��?�m۶m��?      �?      �?              �?      �?        333333�?�������?�������?�������?      �?                      �?      �?        <<<<<<�?�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �Q�٨��?br1���?]��ҟ��?�jc�?      �?        :m��:�?0��b�/�?�u�7[��?Ȥx�L��?      �?        �������?�?              �?GX�i���?�{a���?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?u_[4�?W'u_�?      �?      �?      �?      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?              �?}g���Q�?W�+�ɕ?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?�;�;�?�؉�؉�?_B{	�%�?�^B{	��?B{	�%��?/�����?���Q��?)\���(�?UUUUUU�?UUUUUU�?              �?      �?        (�����?�5��P�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?�������?UUUUUU�?      �?                      �?      �?                      �?�(\����?)\���(�?�������?�������?�Mozӛ�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        �m۶m��?�$I�$I�?333333�?�������?      �?                      �?      �?        333333�?�������?      �?              �?      �?�q�q�?9��8���?      �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?              �?      �?        ��=��?������?�������?�������?              �?      �?        ����^�?^����?UUUUUU�?UUUUUU�?�rv��?�1����?����?�����?X`��??���O?�?�?�������?mЦm�?Y���/Y�?�?<<<<<<�?d!Y�B�?ӛ���7�?�A�A�?��[��[�?              �?      �?      �?�������?�������?      �?                      �?              �?�$I�$I�?�m۶m��?�������?�������?      �?                      �?      �?      �?      �?                      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?'vb'vb�?�a�a�?��y��y�?      �?      �?              �?      �?        (�����?���k(�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�?wwwwww�?      �?                      �?      �?      �?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?      �?              �?      �?                      �?����?����Ǐ�?              �?�?�������?              �?�������?�������?      �?                      �?      �?      �?              �?      �?        �{a���?��=���?�������?�������?      �?      �?              �?      �?                      �?6��P^C�?(������?wwwwww�?�?              �?I�$I�$�?۶m۶m�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ2�3hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKǅ�h��B�1         r                    �?�r,��?�           ��@              e       	          ����?�G�"�?           pz@              <       
             �?(s=u�x�?�            �w@                                  P`@�q�q�?Y             b@                                   �R@�S����?#            �L@                                  �?X�;�^o�?"            �K@                                  0h@և���X�?             @        ������������������������       �                     @        	       
       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�8��8��?             H@                                  @O@���y4F�?             3@                                  �K@�t����?             1@        ������������������������       �                     $@                                   �L@����X�?             @                                  �X@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �                      @               !                    �?�f7�z�?6            �U@                                  �Q@ �Cc}�?             <@        ������������������������       �                      @                                   �g@ ��WV�?             :@                                  `b@      �?             @        ������������������������       �                      @                      	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        "       ;                   xr@TV����?&            �M@       #       ,                    �?ҳ�wY;�?"            �I@        $       %                    X@r�q��?             2@        ������������������������       �                      @        &       '                   �`@�z�G��?             $@        ������������������������       �                     @        (       +                   �d@      �?             @       )       *                    �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        -       :                   Xq@�eP*L��?            �@@       .       /                   `]@���Q��?             9@        ������������������������       �                     @        0       9                    �?      �?             4@       1       2                    �?r�q��?             2@        ������������������������       �                     @        3       4       	          ����?d}h���?
             ,@        ������������������������       �                      @        5       8                   �l@�8��8��?             (@        6       7                    `@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        =       T       	          833�?H�4�l��?�            �m@       >       Q                   �t@ؗp�'ʸ?x            �h@       ?       J                    �?��V�I��?r            �g@        @       I                   �d@r�q��?             >@       A       B                   pb@     ��?
             0@        ������������������������       �                     "@        C       D                    ^@����X�?             @        ������������������������       �                     @        E       F                    �?      �?             @        ������������������������       �                     �?        G       H                     J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             ,@        K       L       	          ����?@=��?_            �c@       ������������������������       �        [            �b@        M       N                     L@؇���X�?             @        ������������������������       �                     @        O       P                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        R       S                     M@      �?              @       ������������������������       �                     @        ������������������������       �                     @        U       V                   `X@�%^�?            �E@        ������������������������       �                     @        W       \                   �j@�����H�?             B@        X       [                   �_@      �?             (@        Y       Z                   `j@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ]       ^                    �? �q�q�?             8@        ������������������������       �                     "@        _       d                   �p@��S�ۿ?
             .@       `       a                    �?؇���X�?             @        ������������������������       �                     @        b       c                     L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        f       k                    @H@z�G�z�?             D@        g       j       	          033@      �?             $@       h       i       
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        l       m                   �c@��S�ۿ?             >@       ������������������������       �                     8@        n       o                    �?�q�q�?             @        ������������������������       �                     @        p       q                    e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        s       �       
             �?l�3/�?�            ps@       t       �                    @G@������?�            �p@        u       �                    �?���N8�?             E@       v       {                    �?�MI8d�?            �B@        w       x       	          833�?X�<ݚ�?             "@        ������������������������       �                      @        y       z                   �a@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        |       }                   �m@@4և���?             <@       ������������������������       �                     1@        ~                          �\@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�����η?�             l@       �       �                    �?�]0��<�?n            �f@       �       �                    �? =[y��?T             a@        ������������������������       �                     4@        �       �                   �_@�8���?E             ]@       �       �                   �[@$�q-�?/            �S@        �       �                    �M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��S�ۿ?-            �R@        �       �                   xt@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                   pl@P�2E��?'            @P@       ������������������������       �                    �C@        �       �                   �Y@ȵHPS!�?             :@        ������������������������       �                     ,@        �       �                    \@      �?
             (@        �       �                   �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     C@        ������������������������       �                    �G@        �       �                    �N@���H��?             E@       �       �                    @M@���B���?             :@       �       �                   Pa@�X�<ݺ?             2@       ������������������������       �                     (@        �       �                   pb@r�q��?             @        �       �                     I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @`@      �?              @       �       �                   �s@�q�q�?             @        ������������������������       �                     @        �       �                   @[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@        �       �                   Xp@d�
��?             F@       �       �                    �?l��
I��?             ;@       �       �                   �k@��s����?             5@       �       �                    b@������?             .@       �       �                   �d@d}h���?
             ,@       �       �                    �?8�Z$���?	             *@        ������������������������       �                     @        �       �                    �M@�<ݚ�?             "@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�t����?
             1@       �       �                   `@�<ݚ�?             "@        ������������������������       �                     @        �       �       	          033�?���Q��?             @       �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  �292ȯ�?�f����?�2t�n��?T�"��?��&:�?���v���?�������?�������?^Cy�5�?(������?J��yJ�?�־a��?۶m۶m�?�$I�$I�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?(������?6��P^C�?�?<<<<<<�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?      �?        O#,�4��?a���{�?%I�$I��?۶m۶m�?              �?O��N���?;�;��?      �?      �?      �?              �?      �?      �?                      �?      �?        u_[4�?E�pR���?�������?�������?UUUUUU�?�������?              �?333333�?ffffff�?              �?      �?      �?      �?      �?              �?      �?                      �?]t�E�?t�E]t�?333333�?�������?              �?      �?      �?�������?UUUUUU�?      �?        I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?              �?      �?        �
j30�?CO��d~�?�S�r
^�?����X�?<�����?AL� &W�?�������?UUUUUU�?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ����&��?�3���y?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?      �?      �?                      �?�}A_��?�}A_�?              �?�q�q�?�q�q�?      �?      �?      �?      �?      �?                      �?      �?        �������?UUUUUU�?      �?        �������?�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ffffff�?ffffff�?      �?      �?�������?UUUUUU�?              �?      �?                      �?�?�������?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?����?;�� y�?B�P�"�?ؽ�u�{�?��y��y�?�a�a�?L�Ϻ��?��L���?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?              �?      �?        �$I�$I�?n۶m۶�?              �?F]t�E�?/�袋.�?      �?                      �?�������?�������?              �?      �?        ������?ų���o�?;ڼOqɠ?\2�h��?�������?�������?              �?a���{�?j��FX�?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?�?�������?�������?�������?              �?      �?        z�z��?_�^��?              �?�؉�؉�?��N��N�?              �?      �?      �?      �?      �?      �?                      �?              �?              �?              �?��y��y�?�0�0�?ى�؉��?��؉���?�q�q�?��8��8�?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�袋.��?�.�袋�?h/�����?Lh/����?�a�a�?z��y���?�?wwwwww�?۶m۶m�?I�$I�$�?;�;��?;�;��?              �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?UUUUUU�?UUUUUU�?              �?      �?        <<<<<<�?�?9��8���?�q�q�?      �?        333333�?�������?      �?      �?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJk�ahG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R��$*     hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK݅�h��B@7         |       
             �?���
%�?�           ��@              m                    �?���Q~�?           �{@              V       	          pff�?�L��d��?�            s@              5                    �?0�� ��?v            �g@                                   �?(옄��?:             W@                      
             �?<ݚ)�?             B@        ������������������������       �                     �?                                  �`@����X�?            �A@       	       
       	          ����?\X��t�?             7@        ������������������������       �                     "@                                   �O@����X�?
             ,@                                 �q@X�<ݚ�?             "@                                  �M@և���X�?             @                     	          ����?      �?             @                                  Pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@               .                    d@h�����?"             L@              +       	          033�?��J�fj�?            �B@                                 @e@�q�q�?             >@                      
             �?z�G�z�?             @        ������������������������       �                     @                                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               *       	          ����?�+e�X�?             9@               !       
             �?����X�?             5@        ������������������������       �                      @        "       %                   �b@���y4F�?             3@        #       $       	          ����?      �?             @        ������������������������       �                     @        ������������������������       �                     @        &       )                    b@$�q-�?             *@       '       (                   l@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ,       -                    N@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        /       0                    �?���y4F�?             3@       ������������������������       �                     &@        1       2                   �m@      �?              @        ������������������������       �                     @        3       4                   �o@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        6       7       	          ����?B�1V���?<            @X@        ������������������������       �                     A@        8       9       	          hff�?���N8�?)            �O@        ������������������������       �                     @        :       I                   P`@z�G�z�?'             N@        ;       D                    �K@`�Q��?             9@       <       C                    @I@r�q��?             2@       =       >                    �?      �?             (@        ������������������������       �                      @        ?       B                   �o@ףp=
�?             $@        @       A       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        E       H                    �?����X�?             @       F       G                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        J       O                    @G@(N:!���?            �A@        K       L       	          033�?�q�q�?             @        ������������������������       �                     �?        M       N                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       S                   �s@      �?             @@       Q       R                   @e@h�����?             <@       ������������������������       �                     ;@        ������������������������       �                     �?        T       U                    w@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        W       j                    `P@�8���?H             ]@       X       [       	          `ff�?��4+̰�?<            @X@        Y       Z                   p@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        \       i                   pp@�x�E~�?6            @V@       ]       b                    �?���U�?$            �L@        ^       _                   �`@      �?             @        ������������������������       �                      @        `       a       	          `ff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        c       d       	          033@�O4R���?!            �J@       ������������������������       �                    �D@        e       h                   �_@�8��8��?             (@        f       g                   �n@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @@        k       l                    �?�S����?             3@        ������������������������       �                     @        ������������������������       �                     0@        n       o                   `Q@г�wY;�?R             a@        ������������������������       �                     �?        p       q                    �?����?�?Q            �`@       ������������������������       �        ?            @Z@        r       w       
             �?ףp=
�?             >@        s       t                    ]@���Q��?             @        ������������������������       �                      @        u       v                    �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        x       y                    @`2U0*��?             9@       ������������������������       �                     2@        z       {                   p@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        }       �       	             �?`>C�#��?�            Pr@       ~       �                    �?�#%�l��?�            �m@              �                    �?���ȑ��?�             j@        �       �       	          @33�?������?             >@       �       �                    �?`�Q��?             9@        �       �                    �L@X�Cc�?	             ,@       ������������������������       �                      @        �       �                   hq@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �g@���!pc�?	             &@        ������������������������       �                     �?        �       �                    ]@z�G�z�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@       �       �                   `l@r�q��?             @        ������������������������       �                     @        �       �                    a@�q�q�?             @        ������������������������       �                     �?        �       �                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @E@P�p�_�?}            `f@        �       �                    ]@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@�E��@�?y            �e@        ������������������������       �        *             N@        �       �                    @��x$�?O            �\@       �       �                    �?������?L             [@       �       �                    @N@hl �&�?C             W@       �       �       	          @33�?���E�??            �U@       ������������������������       �        <            �T@        �       �                   �`@z�G�z�?             @        ������������������������       �                     @        �       �                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   pa@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             0@        ������������������������       �                     @        �       �                    �?������?             ;@        ������������������������       �                      @        �       �                    �?p�ݯ��?             3@       �       �                    �?     ��?             0@        ������������������������       �                     @        �       �                   �b@�	j*D�?	             *@       �       �                    �F@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @K@      �?             @        ������������������������       �                      @        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @b@���b���?$            �L@        �       �                   �b@�������?             >@       �       �                   �Y@8�Z$���?             :@        ������������������������       �                     �?        �       �                    �?H%u��?             9@        ������������������������       �                     �?        �       �                   `]@�8��8��?             8@        ������������������������       �                     @        �       �                   �_@�KM�]�?
             3@        ������������������������       �                     "@        �       �                    �?z�G�z�?             $@        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                   Pa@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�5��?             ;@        ������������������������       �                     $@        �       �                    @ҳ�wY;�?             1@       �       �       	             �?և���X�?
             ,@        ������������������������       �                     @        �       �                    �?���!pc�?	             &@       �       �                    �G@      �?             @        ������������������������       �                      @        �       �                   �e@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��\���?��Q���?ݤ�[r�?���i#�?>��xp�?yp���c�?�4M�4M�?�eY�eY�?ӛ���7�?���,d�?�8��8��?��8��8�?      �?        �$I�$I�?�m۶m��?��Moz��?!Y�B�?              �?�m۶m��?�$I�$I�?r�q��?�q�q�?۶m۶m�?�$I�$I�?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?              �?                      �?n۶m۶�?%I�$I��?к����?�"�u�)�?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?      �?                      �?���Q��?R���Q�?�$I�$I�?�m۶m��?      �?        (������?6��P^C�?      �?      �?              �?      �?        ;�;��?�؉�؉�?UUUUUU�?�������?      �?                      �?              �?              �?۶m۶m�?�$I�$I�?              �?      �?        6��P^C�?(������?      �?              �?      �?              �?�������?�������?      �?                      �?��4l7��?���$2�?              �?��y��y�?�a�a�?      �?        �������?�������?{�G�z�?��(\���?UUUUUU�?�������?      �?      �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        �A�A�?|�W|�W�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?      �?�$I�$I�?�m۶m��?              �?      �?              �?      �?      �?                      �?a���{�?j��FX�? tT����?_\����?      �?      �?      �?                      �?p�\��?����G�?p�}��?	�#����?      �?      �?              �?      �?      �?      �?                      �?�x+�R�?:�&oe�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?^Cy�5�?(������?      �?                      �?�?�?      �?        l�l��?��I��I�?              �?�������?�������?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?{�G�z�?���Q��?              �?�$I�$I�?۶m۶m�?              �?      �?        �$��+6�?7m�AQ'�?4��}yl�?_[4��?��[�)�?�$B�e�?wwwwww�?�?��(\���?{�G�z�?%I�$I��?�m۶m��?      �?        UUUUUU�?�������?      �?                      �?F]t�E�?t�E]t�?              �?�������?�������?              �?�q�q�?�q�q�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        B�D�H�?�7Ck��?      �?      �?      �?              �?      �?              �?      �?        ĦҐs�?E'�卑?      �?        �aܯK*�?��s���?�q�q�?�q�q�?ozӛ���?Y�B��?m��֡�?Ȥx�L��?      �?        �������?�������?      �?              �?      �?      �?                      �?333333�?�������?      �?                      �?      �?              �?        B{	�%��?{	�%���?      �?        ^Cy�5�?Cy�5��?      �?      �?              �?vb'vb'�?;�;��?�q�q�?�q�q�?              �?      �?              �?      �?              �?      �?      �?              �?      �?              �?        1��t��?g1��t�?�������?�������?;�;��?;�;��?      �?        ���Q��?)\���(�?      �?        UUUUUU�?UUUUUU�?              �?(�����?�k(���?              �?�������?�������?              �?�$I�$I�?�m۶m��?�������?333333�?      �?                      �?              �?      �?      �?              �?      �?        h/�����?/�����?      �?        �������?�������?۶m۶m�?�$I�$I�?      �?        t�E]t�?F]t�E�?      �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ6ޤhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�.         h                    �?0����?�           ��@                                  �?������?            |@                      	          ���@�1����?O            ``@                                 �R@`2U0*��?L            @_@        ������������������������       �                     �?                      	             �?�g�y��?K             _@              
                   `X@�T�~~4�?G            @]@               	                    @L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?����X�?D             \@                                   `@���N8�?             5@        ������������������������       �                     $@                                  �`@�C��2(�?	             &@                                  @d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        4            �V@                                   �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               =       
             �?ƹ��"��?�            �s@               &                    �?���N8�?T            `b@                     
             �?��S�ۿ?-            �R@                                  �W@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  pb@����Q8�?*            �Q@       ������������������������       �                     K@                !                     L@������?             1@       ������������������������       �                     &@        "       #                    �M@�q�q�?             @        ������������������������       �                     @        $       %                    �O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        '       0       	          ����?�q�q�?'             R@        (       +                    �?z�G�z�?             9@        )       *                     C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ,       /                   �X@�}�+r��?             3@        -       .                   �W@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        1       <                   8r@JJ����?            �G@       2       5                    �?X��ʑ��?            �E@        3       4                   Pl@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        6       7       
             �?4���C�?            �@@        ������������������������       �                     @        8       9                    �F@l��[B��?             =@        ������������������������       �                     "@        :       ;                    �N@�z�G��?             4@       ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �                     @        >       K       	          ����?�ĚpF�?m            @e@       ?       D                     N@؞�z�̼?L            @]@       @       C                    �?h㱪��?G            �[@        A       B                   `\@���y4F�?
             3@        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �        =            �V@        E       J                    �?և���X�?             @       F       G                    �N@���Q��?             @        ������������������������       �                      @        H       I                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        L       Q                   P`@l`N���?!            �J@        M       P                    �?ףp=
�?             $@        N       O                    �L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        R       S                    �?�^�����?            �E@        ������������������������       �                      @        T       Y                    U@���� �?            �D@        U       X                    c@؇���X�?             @        V       W                    @L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        Z       [                   pi@��hJ,�?             A@        ������������������������       �                     "@        \       ]       	            �?z�G�z�?             9@        ������������������������       �                      @        ^       g                   a@�t����?
             1@        _       `                   �b@�eP*L��?             &@        ������������������������       �                      @        a       f                   �`@�q�q�?             "@       b       e                   �_@؇���X�?             @       c       d                   �j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        i       t                    �?��8���?�            �q@        j       o       	          ����?j���� �?             A@        k       l                     N@�8��8��?             (@       ������������������������       �                      @        m       n       	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        p       q       	          ����?��2(&�?             6@       ������������������������       �        
             .@        r       s                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        u       �                    @G@|�(��?�            �o@        v       }                    @F@     ��?             @@       w       x       	          ����?�C��2(�?             6@        ������������������������       �                     $@        y       |                   �l@r�q��?             (@        z       {                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ~                          @`@      �?             $@        ������������������������       �                      @        �       �                   �Z@      �?              @        ������������������������       �                     @        �       �                   �k@���Q��?             @        ������������������������       �                      @        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?�L�3�?�            �k@       �       �                    a@����$}�?z            @g@       �       �                   i@`'�J�?d             c@        ������������������������       �        '             N@        �       �                   �\@`Jj��?=            @W@        ������������������������       �                     @        �       �                    �R@(;L]n�?;            �V@       �       �                   �[@�D�e���?9            @U@        �       �                     P@�FVQ&�?            �@@       �       �                    �O@�8��8��?             8@       �       �                   `[@P���Q�?             4@       ������������������������       �                     2@        �       �                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          :33�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �        %             J@        �       �                   �b@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   0a@6YE�t�?            �@@        ������������������������       �                      @        �       �                    @��a�n`�?             ?@       �       �       	          ����?��S�ۿ?             >@        ������������������������       �                     $@        �       �                   �[@ףp=
�?             4@        ������������������������       �                     �?        �       �                    q@�}�+r��?             3@       ������������������������       �                     &@        �       �                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �d@������?             A@       �       �                   �a@     ��?             @@       �       �                   �`@�8��8��?             8@        ������������������������       �                     (@        �       �                    �?r�q��?             (@       �       �                   Pa@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                   @\@z�G�z�?             @        ������������������������       �                     @        �       �                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ���^L�?���Y�?I�$I�$�?n۶m۶�?J�eDP�?����?���Q��?{�G�z�?              �?��{���?�B!��??�s?�s�?���?�������?�������?      �?                      �?n۶m۶�?�$I�$I�?��y��y�?�a�a�?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?              �?      �?                      �?��`=��?�P�?�w�?��y��y�?�a�a�?�?�������?      �?      �?      �?                      �?��Vج?O�o�z2�?              �?�?xxxxxx�?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        (�����?�5��P�?�������?�������?              �?      �?                      �?��
br�?x6�;��?��}A�?�}A_�?�������?�������?      �?                      �?m��&�l�?'�l��&�?      �?        ���=��?GX�i���?      �?        333333�?ffffff�?              �?      �?              �?        �������?�������?^�^��?�ꡮ?־a���?��)A��?6��P^C�?(������?              �?      �?              �?        �$I�$I�?۶m۶m�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �R���?
�[���?�������?�������?�������?�������?              �?      �?                      �?�5eMYS�?֔5eMY�?              �?jW�v%j�?,Q��+�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?KKKKKK�?�������?      �?        �������?�������?      �?        �������?�������?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �L[����?�,)D��?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        t�E]t�?��.���?              �?۶m۶m�?�$I�$I�?              �?      �?        ��i��i�?-˲,˲�?      �?      �?F]t�E�?]t�E�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?־a��?=%�S�<�?Hy�G�?n���?�?�������?              �?�B!��?���{��?      �?        �?�������?�???????�?|���?>����?UUUUUU�?UUUUUU�?�������?ffffff�?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?              �?              �?�������?�������?              �?      �?        e�M6�d�?'�l��&�?      �?        �c�1Ƹ?�s�9��?�?�������?              �?�������?�������?      �?        (�����?�5��P�?              �?      �?      �?      �?                      �?      �?        �?xxxxxx�?      �?      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?F]t�E�?]t�E�?      �?                      �?      �?              �?      �?�������?�������?              �?      �?      �?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��{hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�-         f                    �?�ܲ�}��?�           ��@              ;       
             �?��B��?�            Pz@              6                    c@�M�u�?�            �s@                                 Pe@��L~1_�?�            0p@        ������������������������       �        (             P@               1                    �?z�G�z�?q            `h@                                 �e@�<ݚ�?_            `e@        ������������������������       �                     @        	       0                   �a@��%c�?^            �d@       
       %       	             �?T�iA�?O            �a@                                   �?���`��?             �P@                                   `@r�q��?             2@        ������������������������       �                     "@                                   �?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @                                  �[@�J��%�?            �H@                                   �N@X�Cc�?             ,@                                 �`@      �?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               $                   �e@z�G�z�?            �A@              #                    @M@      �?             @@                     	          ����?�㙢�c�?             7@        ������������������������       �                     "@                                   �?����X�?	             ,@        ������������������������       �                     @               "                   �s@      �?              @                     	          hff�?�q�q�?             @        ������������������������       �                     �?                !                   �m@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        &       +                   `i@��pBI�?/            @R@        '       (                    �?z�G�z�?             @        ������������������������       �                      @        )       *                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ,       -                   0c@ ��ʻ��?,             Q@       ������������������������       �        *            �P@        .       /                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        2       5       
             �? �q�q�?             8@        3       4                   `v@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        7       8                    `R@ �Jj�G�?!            �K@       ������������������������       �                    �I@        9       :       	             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        <       G                   @E@�"��61�?E            �Z@        =       D                   @b@؇���X�?             5@       >       C                   @^@      �?             0@        ?       @                    �?z�G�z�?             @        ������������������������       �                      @        A       B       	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        E       F                    d@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        H       ]                    �?2X��ʑ�?6            �U@       I       T                    �L@     ��?)             P@       J       S                    �?=QcG��?             �G@        K       L                   0n@      �?             (@        ������������������������       �                     @        M       N                   po@      �?              @        ������������������������       �                      @        O       R                   `\@r�q��?             @        P       Q                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �A@        U       Z                   �l@��.k���?	             1@       V       W                    a@�<ݚ�?             "@       ������������������������       �                     @        X       Y                   @c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        [       \                   �e@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ^       e       	          ����?�X����?             6@       _       `                    �?      �?             ,@        ������������������������       �                     @        a       d                   �p@���|���?             &@        b       c                    @K@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        g       �                    �?�,�;i��?�            �s@       h       �       	          033�?>�<���?�            �p@       i       j                   `R@d���A�?�             n@        ������������������������       �                     @        k       p                    �?hV'���?�            `m@        l       o                    �? qP��B�?6            �U@        m       n                    �?�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �        .            �Q@        q       v                   �h@�3�o���?X            �b@        r       u                    �?`���i��?             F@        s       t                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     E@        w       �                     L@4�2%ޑ�?A            @Z@       x       }                     B@      �?-             R@        y       |                   @p@�z�G��?             $@        z       {       
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ~       �       
             �?��a�n`�?(             O@               �                   f@�eP*L��?             &@       �       �                   �o@      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �I@        �       �                    �Q@�eP*L��?            �@@       �       �                   �Z@���Q��?             >@        ������������������������       �                     @        �       �                    �L@      �?             8@        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                   Hp@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          pff�?      �?             0@       ������������������������       �                     &@        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                   �c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �? �o_��?             9@       �       �                    �?؇���X�?             5@       �       �                   @a@���!pc�?             &@        ������������������������       �                     �?        �       �       
             �?z�G�z�?             $@       �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                    �N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                   �i@��|�5��?!            �G@        �       �                   �e@�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?        �       �       	          `ff�?J�8���?             =@       �       �                   �j@��X��?             <@        ������������������������       �                      @        �       �       	          ����?R�}e�.�?             :@       �       �       
             �?�q�q�?             5@       �       �                   �`@�<ݚ�?             2@       ������������������������       �                     &@        �       �                   m@և���X�?             @        ������������������������       �                     @        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  ����u��?/�E��?s�XV
�?#�ij=?�?�n�{DN�?H��n��?c4�w-F�?��t.�?              �?�������?�������?�q�q�?9��8���?      �?        GS��r�?.+Jx��?��+��+�?PuPu�?�1����?*g��1�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?9/����?c}h���?%I�$I��?�m۶m��?      �?      �?              �?      �?              �?        �������?�������?      �?      �?d!Y�B�?�7��Mo�?              �?�$I�$I�?�m۶m��?              �?      �?      �?UUUUUU�?UUUUUU�?      �?        333333�?�������?              �?      �?                      �?              �?      �?        ����?���Ǐ�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�������?              �?      �?      �?              �?      �?                      �?UUUUUU�?�������?      �?      �?              �?      �?                      �?��)A��?k߰�k�?              �?      �?      �?              �?      �?        9��/Ċ�?��L�w��?�$I�$I�?۶m۶m�?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?333333�?      �?                      �?}A_���?}A_��?      �?      �?x6�;��?AL� &W�?      �?      �?      �?              �?      �?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �?�������?9��8���?�q�q�?      �?              �?      �?              �?      �?              �?      �?              �?      �?        ]t�E]�?�E]t��?      �?      �?              �?]t�E]�?F]t�E�?�������?�������?              �?      �?              �?                      �?F܋��?u�G���?֝VwZ��?���"���?F�F��?�熑��?              �?����R�?�"��i�?��}A�?�}A_З?�������?�?      �?                      �?      �?        �a�ۀ��?ExR��y�?F]t�E�?F]t�E�?      �?      �?              �?      �?              �?        �������?�A�A�?      �?      �?ffffff�?333333�?      �?      �?              �?      �?              �?        �s�9��?�c�1Ƹ?]t�E�?t�E]t�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        t�E]t�?]t�E�?333333�?�������?              �?      �?      �?      �?      �?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?      �?        333333�?�������?              �?      �?      �?      �?                      �?              �?�Q����?
ףp=
�?�$I�$I�?۶m۶m�?t�E]t�?F]t�E�?      �?        �������?�������?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        x6�;��?br1���?�q�q�?��8��8�?              �?      �?        |a���?�rO#,��?%I�$I��?n۶m۶�?      �?        �;�;�?'vb'vb�?UUUUUU�?UUUUUU�?�q�q�?9��8���?              �?�$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ?{�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKͅ�h��B@3         �       
             �?8}�ý�?�           ��@              _                   �b@�B�@�L�?           �z@              6                   P`@`����e�?�            �v@                                  �?`.��A��?�            �m@                                   i@�q�q�?             2@                      	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        	                           `P@d}h���?             ,@       
                          ps@�8��8��?	             (@       ������������������������       �                     $@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                  �Q@��Au5a�?�            �k@                      
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                      	             �?�2����?�            `k@        ������������������������       �                     �J@               +                    �?���Ehz�?i            �d@                     	          ����?Xl���?I            �\@        ������������������������       �                     @                                  �[@�v�ɱ?H            �[@        ������������������������       �                     G@               *                    �Q@����?,            @P@              !                    �D@�i�y�?*            �O@                                   b@      �?              @       ������������������������       �                     @                                    �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        "       #                    @L@ �Jj�G�?$            �K@       ������������������������       �                    �@@        $       )                    �L@���7�?             6@        %       &                   �d@z�G�z�?             @        ������������������������       �                      @        '       (                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                      @        ,       5                   p`@ȵHPS!�?              J@        -       4                   �^@�z�G��?             4@       .       /                   �^@���Q��?	             .@        ������������������������       �                     @        0       1       
             �?      �?             (@        ������������������������       �                      @        2       3                    �L@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @@        7       P                    �?�<jV�?J            �^@        8       ?                   �h@F�����?            �F@        9       :                   0a@���N8�?             5@        ������������������������       �                     (@        ;       >                    b@�����H�?             "@        <       =                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        @       G                    �K@�q�q�?             8@        A       B                   �\@"pc�
�?             &@        ������������������������       �                     �?        C       F       	          @33�?ףp=
�?             $@        D       E                   �a@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        H       I                   p`@��
ц��?	             *@        ������������������������       �                     @        J       O       	           33@�q�q�?             "@       K       L                   0b@؇���X�?             @       ������������������������       �                     @        M       N                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        Q       X                    �?ȵHPS!�?-            �S@       R       W                    �G@�U�=���?&            �P@        S       T                     F@�E��ӭ�?	             2@       ������������������������       �                     (@        U       V       	             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     H@        Y       Z                   �a@�q�q�?             (@        ������������������������       �                     @        [       \                    �?�����H�?             "@        ������������������������       �                     @        ]       ^                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        `       a                    �A@$/����?+            @P@        ������������������������       �                     @        b       k       	          ����?�^�����?)             O@        c       d                    c@�<ݚ�?             2@        ������������������������       �                      @        e       j                    �?      �?
             0@       f       i                    �?"pc�
�?             &@        g       h                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        l                           �?�X���?             F@       m       v                    �?4�2%ޑ�?            �A@        n       q                   0p@      �?             0@        o       p       	          033�?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        r       s                    �?      �?              @        ������������������������       �                     @        t       u                    @N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        w       ~                   0m@�KM�]�?             3@       x       }                   �l@z�G�z�?             $@       y       z                   @e@�����H�?             "@       ������������������������       �                     @        {       |                    �I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �       
             �?�<ݚ�?             "@        ������������������������       �                     �?        �       �       	          433�?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ���@�Ƒ�*�?�            0s@       �       �                    �?H;T*St�?�            `r@        �       �       	          ����?z�J�?A            �W@       �       �                    �?z�G�z�?/            @P@       �       �                    �I@���*�?*             N@        �       �                    �?      �?             @@        �       �                   �c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        �       �                    @J@X�Cc�?             <@        ������������������������       �                      @        �       �                   e@�	j*D�?             :@       �       �                    `@ �o_��?             9@        �       �                    �K@r�q��?	             (@        ������������������������       �                     �?        �       �                   d@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                    @N@�n_Y�K�?	             *@       �       �                    b@z�G�z�?             $@        ������������������������       �                     @        �       �                     M@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          833�?���Q��?             @       �       �                     L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    @E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    b@����"�?             =@       �       �                   �Y@���y4F�?             3@        ������������������������       �                      @        �       �                    �?�t����?
             1@        ������������������������       �                     �?        �       �                    �?      �?	             0@       �       �       	          ����?�����H�?             "@       ������������������������       �                     @        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �c@�z�G��?             $@       �       �       	          ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       	            �?`2U0*��?}             i@       �       �                    �O@@���I�?b            �c@       ������������������������       �        \            `b@        �       �                   Pc@ףp=
�?             $@       ������������������������       �                      @        �       �                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �_@�T|n�q�?            �E@        �       �                     L@�q�q�?             (@       �       �                    �I@r�q��?             @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ?@        ������������������������       �                     *@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  a[ӿc�?PR Np�?��v��?�@�Rb�?X�s��C�?jc��?@|4!/l�?xp�zR�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?        ۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        �7�7�?�����?      �?      �?      �?                      �?H�!��d�?��m���?              �?���\V�?A	o4u~�?��Gp�?��>���?      �?        5'��Ps�?��w����?              �? �����?~�~��?AA�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ��)A��?k߰�k�?              �?F]t�E�?�.�袋�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �؉�؉�?��N��N�?333333�?ffffff�?�������?333333�?              �?      �?      �?      �?        �������?333333�?      �?                      �?              �?              �?鰑�?<�œ[<�?؂-؂-�?�>�>��?�a�a�?��y��y�?              �?�q�q�?�q�q�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?/�袋.�?F]t�E�?              �?�������?�������?�������?�������?      �?                      �?      �?        �;�;�?�؉�؉�?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?        �؉�؉�?��N��N�?e�M6�d�?�M6�d��?r�q��?�q�q�?              �?�������?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?              �?�������?�������?      �?                      �?�?�?�? �����?              �?!�B�?���{��?�q�q�?9��8���?      �?              �?      �?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?]t�E�?�E]t��?�������?�A�A�?      �?      �?      �?      �?      �?                      �?      �?      �?              �?      �?      �?      �?                      �?�k(���?(�����?�������?�������?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �q�q�?9��8���?      �?              �?      �?      �?                      �?dXn��?�o��G��?�r
^N��??4և���?��
br�?�w6�;�?�������?�������?""""""�?wwwwww�?      �?      �?�������?�������?              �?      �?              �?        %I�$I��?�m۶m��?              �?vb'vb'�?;�;��?
ףp=
�?�Q����?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?                      �?;�;��?ى�؉��?�������?�������?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        �i��F�?	�=����?(������?6��P^C�?      �?        �?<<<<<<�?      �?              �?      �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?ffffff�?333333�?۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���Q��?{�G�z�?jX���?Kz��z?      �?        �������?�������?      �?              �?      �?              �?      �?        ���)k��?6eMYS��?�������?�������?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��}whG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@,         f       
             �?\\��?�           ��@              A                   �a@���;�?	           @{@                                  �?$�q-�?�            �s@                                  �a@؇���X�?1             U@                                 @R@d}h���?"             L@        ������������������������       �                     @                                  �X@8�Z$���?!             J@                                    M@�q�q�?             "@        	       
       	             ���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?X�EQ]N�?            �E@                                  @O@r�q��?             >@                                  �? �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@                      	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     <@                      
             �?�}�+r��?�            �l@                                  �r@      �?             @@       ������������������������       �                     =@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               8                   �_@�ib�=�?|            �h@              5       	          ���@ 	��p�?Z             b@                                   @L@���?S            �`@        ������������������������       �        %             N@        !       4       	          ����?H0sE�d�?.            �R@       "       '                    �L@PN��T'�?!             K@        #       $                   @_@և���X�?             @        ������������������������       �                     @        %       &                   �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        (       3                   �`@dP-���?            �G@        )       .                    _@���|���?             &@       *       +                    �?r�q��?             @       ������������������������       �                     @        ,       -       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        /       0                    [@���Q��?             @        ������������������������       �                      @        1       2                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     B@        ������������������������       �                     5@        6       7                   �_@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        9       :                   �m@���J��?"            �I@       ������������������������       �                    �A@        ;       @       	          ����?      �?             0@        <       =                    �?�q�q�?             @        ������������������������       �                     �?        >       ?                   ps@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             *@        B       C                   �h@0�n�"��?H             _@        ������������������������       �                     8@        D       U                   pn@x��#���?:             Y@        E       J                    �K@�D��?            �H@       F       I                   �\@`Jj��?             ?@        G       H       	          ����?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     8@        K       N                   b@b�2�tk�?
             2@        L       M                    �L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        O       P                    @M@�θ�?             *@        ������������������������       �                     @        Q       T                    @P@      �?             @       R       S                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        V       e                    f@�t����?            �I@       W       X                   �b@z�G�z�?            �F@        ������������������������       �                     &@        Y       Z                     J@�������?             A@        ������������������������       �                     ,@        [       `                    �?�G�z��?             4@        \       ]                    �K@z�G�z�?             $@        ������������������������       �                     @        ^       _                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        a       b       	          `ff�?ףp=
�?             $@       ������������������������       �                     @        c       d                     M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        g       �                    �?��P�;�?�            �r@       h       s                    �?����!�?�            �n@        i       l                    @C@X��%�?5            �U@        j       k                    �?���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        m       n                   Pt@�e���@�?0            @S@       ������������������������       �        ,            �Q@        o       p                     M@r�q��?             @        ������������������������       �                     @        q       r                    �O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        t       �                    �?l������?g            �c@        u       x                   @E@ҳ�wY;�?            �I@        v       w       	          ����?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        y       z                   �b@:�&���?            �C@        ������������������������       �                     1@        {       |                   �i@�X����?             6@        ������������������������       �                     @        }       �                     L@�t����?             1@       ~       �                   `\@��S�ۿ?
             .@               �                    �E@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �L@�F�1G�?H            �Z@       �       �       	             @����ȫ�?<            �T@       ������������������������       �        ;            @T@        ������������������������       �                     �?        �       �                   `l@���Q��?             9@        �       �       	            �?r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �       	             �?�n_Y�K�?             *@       �       �       	          @33�?���!pc�?             &@       �       �                   @c@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �K@Fmq��?            �J@        �       �                    �?���!pc�?	             &@       �       �                     J@���Q��?             @       �       �                   pj@      �?             @        ������������������������       �                      @        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?��i#[�?             E@        �       �                    �Q@�q�q�?             (@       �       �                   �f@�<ݚ�?             "@       �       �                    h@      �?              @        �       �                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?             >@        ������������������������       �                     �?        �       �                   q@д>��C�?             =@       �       �                   �`@؇���X�?             <@       ������������������������       �                     0@        �       �                   �`@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B  �+�U�?�js��?K`�~��?�'K`�~�?;�;��?�؉�؉�?�$I�$I�?۶m۶m�?۶m۶m�?I�$I�$�?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?                      �?qG�wĽ?w�qG�?UUUUUU�?�������?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?(�����?�5��P�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        /�����?����>4�?�{a���?������?t��:W�?��oS��?              �?O贁N�?��b�/��?h/�����?&���^B�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?        W�+�ɵ?�����F�?F]t�E�?]t�E]�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�������?      �?                      �?�?______�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?SJ)��R�?�Zk����?              �?R���Q�?\���(\�?������??4և���?���{��?�B!��?�m۶m��?�$I�$I�?              �?      �?              �?        9��8���?�8��8��?�������?�������?              �?      �?        �؉�؉�?ى�؉��?              �?      �?      �?      �?      �?              �?      �?                      �?�������?�������?�������?�������?              �?�������?�������?              �?�������?�������?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �{��6`�?.�$�?�����?K��o!`�? ��2)�?��֡�l�?333333�?�������?              �?      �?        qV~B���?�cj`?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        :�g *�?7a~W��?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?�A�A�?�o��o��?      �?        �E]t��?]t�E]�?              �?<<<<<<�?�?�������?�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?�;u-7�?�+J�#�?������?������?      �?                      �?�������?333333�?UUUUUU�?�������?      �?                      �?;�;��?ى�؉��?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?                      �?      �?                      �?~�	�[�?�x+�R�?F]t�E�?t�E]t�?�������?333333�?      �?      �?              �?      �?      �?      �?                      �?      �?              �?        �<��<��?�a�a�?�������?�������?9��8���?�q�q�?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?�������?�������?      �?        |a���?a���{�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�,�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�-         V       	          ����?.��X~��?�           ��@              -                    �?�S
�T�?�            �w@                      
             �?�99lMt�?b            �c@              	                    �?�Ra����?8             V@                                   �?      �?             @        ������������������������       �                      @                      	          @33�?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        
              	          833�?ĴF���?2            �T@       ������������������������       �        (            �Q@                                   b@�q�q�?
             (@                                  �I@�z�G��?             $@        ������������������������       �                      @                                   _@      �?              @                                  �\@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @               ,                   0e@�!���?*             Q@              +                   �f@��Q:��?$            �M@                                 @E@���dQ'�?#            �L@                      	          ����?d}h���?	             ,@                                  �]@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               &                    @M@RB)��.�?            �E@              !                     E@��S�ۿ?             >@                                   �[@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        "       %                    ]@`2U0*��?             9@        #       $                    �I@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        '       *                     P@��
ц��?             *@       (       )                   �a@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        .       G       
             �?���,��?�            �k@        /       6                   �c@�s��:��?             C@        0       1                    V@�����H�?             "@        ������������������������       �                     @        2       5                    @z�G�z�?             @       3       4                   `X@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        7       F       	          833�?П[;U��?             =@       8       E                    �?\X��t�?             7@       9       @                    �?�\��N��?             3@        :       ?       	          ����?z�G�z�?             $@       ;       >                   �o@      �?              @       <       =                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        A       D                   �`@�<ݚ�?             "@        B       C                   @\@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        H       O                   �s@��<b�ƥ?q             g@       I       J                    @L@@c����?i            @e@       ������������������������       �        [            �b@        K       N                    �L@���7�?             6@        L       M                    c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@        P       Q                   �`@d}h���?             ,@       ������������������������       �                     "@        R       S                   0c@���Q��?             @        ������������������������       �                      @        T       U                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        W       �                    �?2�x���?�            @v@        X       w       	          033�?J!�k���?M             `@       Y       l                   �b@      �?/             T@       Z       k                   r@Hث3���?            �C@       [       \                   `\@      �?             @@        ������������������������       �                     @        ]       j                    �?�q�����?             9@       ^       e                   �a@�q�q�?             2@       _       d                    �?"pc�
�?             &@       `       c       	             �?���Q��?             @       a       b                    �M@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        f       i                    �?և���X�?             @        g       h                    �K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        m       v                   Pm@���?            �D@        n       u                    �?�G��l��?             5@       o       p                   Pc@j���� �?	             1@        ������������������������       �                     @        q       t       	          ����?����X�?             ,@       r       s                   �f@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     4@        x       �                    �? \� ���?            �H@        y       �                   d@H%u��?             9@       z       {                   `c@�8��8��?             8@       ������������������������       �        
             1@        |       }                   `Z@����X�?             @        ������������������������       �                     @        ~                           �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   ``@      �?             8@       �       �       	          ��� @�q�q�?	             (@       �       �                     H@      �?              @        ������������������������       �                     @        �       �                   @_@�q�q�?             @       �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �       	          ����?�C&�l��?�            `l@        �       �                   �c@t����?B            �Z@       �       �                     F@p���p�?A            �Y@        �       �                   �\@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          033�?p�qG�?=             X@       �       �                    �?Pa�	�?)            �P@       ������������������������       �                      J@        �       �                   �_@؇���X�?	             ,@       ������������������������       �                     $@        �       �                   @k@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @L@ףp=
�?             >@       ������������������������       �                     6@        �       �                    �M@      �?              @        �       �       
             �?      �?             @       �       �                    ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �Z@Xsj�]�?R            @^@        ������������������������       �                     �?        �       �                    @�(\����?Q             ^@       �       �                    �? ����?P            �]@       �       �       	          ��� @`�߻�ɒ?G             [@       �       �                    �M@ pƵHP�?$             J@       ������������������������       �                     @@        �       �                   �`@P���Q�?             4@       ������������������������       �                     (@        �       �                    Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        #             L@        �       �                    �?�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  ��� ���?���o���?�V�Zk�?�RJ�)�?�o��o��?5H�4H��?]t�E�?]t�E]�?      �?      �?      �?              �?      �?              �?      �?        ە�]�ڵ?E�JԮD�?              �?�������?�������?ffffff�?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?�������?'u_[�?�A�I��?ZLg1���?Lg1��t�?۶m۶m�?I�$I�$�?۶m۶m�?�$I�$I�?      �?                      �?              �?S֔5eM�?���)k��?�������?�?�������?�������?              �?      �?        ���Q��?{�G�z�?�������?UUUUUU�?      �?                      �?      �?        �؉�؉�?�;�;�?t�E]t�?]t�E�?      �?                      �?              �?              �?      �?        X��;ze�?C�I .Լ?�k(���?��k(��?�q�q�?�q�q�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�{a���?��=���?��Moz��?!Y�B�?y�5���?�5��P�?�������?�������?      �?      �?      �?      �?              �?      �?              �?              �?        �q�q�?9��8���?�������?333333�?              �?      �?                      �?              �?      �?        ��7��M�?d!Y�B�?�������?x?      �?        �.�袋�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        I�$I�$�?۶m۶m�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        �3��g�?s����?�'�	{��?(�	{�?      �?      �?��-��-�?�i�i�?      �?      �?              �?���Q��?�p=
ף�?UUUUUU�?UUUUUU�?/�袋.�?F]t�E�?333333�?�������?      �?      �?      �?                      �?      �?              �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?              �?      �?        28��1�?8��18�?1�0��?��y��y�?ZZZZZZ�?�������?      �?        �$I�$I�?�m۶m��?F]t�E�?]t�E�?              �?      �?              �?              �?              �?        և���X�?
^N��)�?���Q��?)\���(�?UUUUUU�?UUUUUU�?              �?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?              �?              �?      �?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?UUUUUU�?�������?      �?                      �?�<.}�+�?c8Z����?:�&oe�?y+�R�?C��ڸ?�E|���?�m۶m��?�$I�$I�?              �?      �?        �������?UUUUUU�?|���?|���?              �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �������?�������?              �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?        ���k��?7�A�0��?      �?        �������?333333�?�5�5�?�Qv�Qv�?h/�����?B{	�%��?;�;��?'vb'vb�?              �?�������?ffffff�?              �?      �?      �?      �?                      �?              �?F]t�E�?]t�E�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�%\hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKم�h��B@6         `       	          ����?�_y���?�           ��@              +                    �?b���L��?�            @x@                                   �?l�;�	�?Z            �b@                                 �Y@��V�I��?;            �W@        ������������������������       �                     @                                  �_@ƈ�VM�?9            @V@                                  �Z@���}<S�?             7@        ������������������������       �                     &@        	       
                    [@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@                      
             �?r٣����?,            �P@                                  0i@ҳ�wY;�?
             1@                                  �_@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                                  �b@ i���t�?"            �H@       ������������������������       �                     9@                                   �M@�q�q�?             8@                                 `\@ףp=
�?             4@                                   q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@                                   a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               *                   `c@�>4և��?             L@              #                   ``@�d�����?             C@                                  q@���N8�?             5@       ������������������������       �                     3@        !       "                   Pa@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       '       
             �?��.k���?
             1@        %       &       	             �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        (       )       	             �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     2@        ,       I       
             �?�p�I�?�            �m@        -       4                    �?J�8���?$             M@        .       3       	          ����?     ��?             0@       /       0                    �I@�n_Y�K�?             *@        ������������������������       �                     @        1       2                     P@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        5       H                    �?d}h���?             E@       6       A       	          ����?$��m��?             :@       7       @                    �L@���y4F�?             3@       8       ?                   o@���|���?	             &@       9       >                    �?      �?              @       :       =                    �?�q�q�?             @       ;       <                   0a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        B       G                    �N@����X�?             @       C       F                    �?���Q��?             @       D       E                    @L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        J       Y                    �?(;L]n�?e            �f@       K       R                   pa@������?[            `d@       L       M       	            �? 4^��?C            �]@       ������������������������       �        >            �[@        N       O                    �?�����H�?             "@        ������������������������       �                     @        P       Q                   �_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        S       T                    �N@t��ճC�?             F@       ������������������������       �                    �B@        U       V                   Pb@և���X�?             @        ������������������������       �                     @        W       X                    s@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       _                    �?�t����?
             1@        [       ^                    �?���Q��?             @        \       ]                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        a       �                   �b@2�8XF��?�            �u@       b       �                    �?p���A�?�             r@       c       �       
             �?��^ҺR�?�            �l@       d       g       	          ����?�����?�            �h@        e       f                   @e@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        h       �                    �Q@p�q��?~             h@       i       ~                   {@��R�x��?{            `g@       j       w       	          033@�:�5ӣ�?y             g@       k       p                    �?@��t��?`             b@        l       o                   @_@8�Z$���?	             *@        m       n                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        q       v                    @G@�\5ݓˎ?W            �`@        r       s                    �?��S�ۿ?             .@       ������������������������       �        
             *@        t       u                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        K            @]@        x       }                    �J@ףp=
�?             D@        y       z                   pk@և���X�?             @        ������������������������       �                      @        {       |                    @J@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �@@               �                   ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �_@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    c@      �?             @@       �       �                   �u@H%u��?             9@       �       �                   �^@�8��8��?             8@        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                    @M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             2@        ������������������������       �                     �?        �       �       	             �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �_@L
�q��?(            �M@       �       �                    @"pc�
�?            �@@       �       �                    �?�r����?             >@        �       �                    �P@���!pc�?             &@       �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          033�?�q�q�?             @        ������������������������       �                     �?        �       �                    @R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�}�+r��?             3@       �       �                   P`@�C��2(�?             &@        �       �                   �\@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   Xq@��
ц��?             :@       �       �                   �c@���|���?             6@       �       �                    �?��.k���?             1@       �       �       	          ����?�q�q�?             (@        �       �                   �a@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                   @a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @N@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @L@l��[B��?%             M@       �       �                    �?�������?             A@        �       �       	          `ff�?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �[@`�Q��?             9@        ������������������������       �                     @        �       �                    �C@��s����?             5@        �       �                    �B@      �?             @       �       �                   �r@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�t����?	             1@       ������������������������       �                     &@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?�q�q�?             8@        �       �                    �?      �?             @       �       �                    �M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   c@�����H�?             2@        ������������������������       �                     �?        �       �                    �?�IєX�?             1@       ������������������������       �                     &@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  V�.�#��?աh6n��?����?�:*���?t�@�t�?ƒ_,���?G}g����?r1����?              �?+Y�JV��?�MmjS��?d!Y�B�?ӛ���7�?              �?UUUUUU�?�������?      �?                      �?>���>�?|���?�������?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?/�����?����X�?      �?        UUUUUU�?�������?�������?�������?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?�m۶m��?�$I�$I�?y�5���?Cy�5��?�a�a�?��y��y�?              �?      �?      �?      �?                      �?�������?�?�$I�$I�?۶m۶m�?              �?      �?        �������?�������?      �?                      �?              �?:�:��?���?|a���?�rO#,��?      �?      �?;�;��?ى�؉��?      �?        �$I�$I�?�m۶m��?              �?      �?              �?        ۶m۶m�?I�$I�$�?vb'vb'�?�N��N��?(������?6��P^C�?F]t�E�?]t�E]�?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?              �?              �?              �?�m۶m��?�$I�$I�?333333�?�������?      �?      �?      �?                      �?              �?      �?                      �?�������?�?�x�%�6�?)��I� �?�(��(��?�5�5�?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?        �E]t��?t�E]t�?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?<<<<<<�?�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ����D�?V����n�?��8��8�?�q�q�?����y�?��G���?�����?/,FBi��?�������?333333�?              �?      �?        UUUUUU�?�����*�?�и[�?��rD���?�5!({_�?��}M��?��RA�/�?*h���V�?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?              �?|��?�|���?�?�������?              �?      �?      �?              �?      �?                      �?�������?�������?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?                      �?      �?      �?      �?                      �?333333�?�������?      �?                      �?      �?      �?���Q��?)\���(�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �m۶m��?�$I�$I�?              �?      �?        �pR���?��V'�?F]t�E�?/�袋.�?�?�������?t�E]t�?F]t�E�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?(�����?�5��P�?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �;�;�?�؉�؉�?]t�E]�?F]t�E�?�������?�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?�������?333333�?      �?              �?      �?      �?                      �?�������?�������?              �?      �?              �?                      �?���=��?GX�i���?�������?�������?�q�q�?�q�q�?              �?      �?        ��(\���?{�G�z�?              �?z��y���?�a�a�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?<<<<<<�?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?      �?      �?      �?              �?      �?                      �?�q�q�?�q�q�?      �?        �?�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ2�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@=         �                    �?~�w�H�?�           ��@              �                    @N@BA�V�?           �{@              :                   P`@>���b�?�            pt@              1       
             �?�:�B��?j             f@                     	             �?������?W            @b@        ������������������������       �                     =@                                  �R@�����H�?D            @]@        ������������������������       �                     @        	                           �?x�}b~|�?C            �\@        
                            L@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @                                  �_@�q-�?=             Z@                                  �^@\-��p�?             =@                                  k@���}<S�?             7@                                  `_@      �?              @        ������������������������       �                     @                                   �?���Q��?             @                      	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@                                  @]@�q�q�?             @                                  �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               0                   �b@`2U0*��?,            �R@                                  �D@�}�+r��?#            �L@        ������������������������       �                     �?                !                    @K@h�����?"             L@        ������������������������       �                     8@        "       /                   �a@      �?             @@       #       $       
             �?���}<S�?             7@        ������������������������       �                      @        %       &                    �?�����?             5@        ������������������������       �                     @        '       (                   �X@�����H�?             2@        ������������������������       �                     �?        )       .                    �?�IєX�?
             1@       *       +                   �j@؇���X�?             @       ������������������������       �                     @        ,       -                   �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     "@        ������������������������       �        	             2@        2       3       	          ����?`՟�G��?             ?@       ������������������������       �        
             .@        4       5                    �?      �?	             0@        ������������������������       �                     �?        6       7                    �M@��S�ۿ?             .@       ������������������������       �                     $@        8       9                   �]@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ;       d                    �?*;L]n�?]            �b@       <       ?                    @C@~�hP��?0            �R@        =       >                   `]@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        @       M       
             �?:-�.A�?+            �P@        A       L                    �?���Q��?             4@       B       C                    a@և���X�?	             ,@        ������������������������       �                     @        D       G                    �F@�q�q�?             "@        E       F                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        H       I                   �`@r�q��?             @       ������������������������       �                     @        J       K       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        N       c                    �?��0{9�?            �G@       O       Z                    �?��r._�?            �D@        P       W                   d@�t����?             1@       Q       R                    q@@4և���?             ,@        ������������������������       �                     "@        S       V                    �?z�G�z�?             @       T       U                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        X       Y                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        [       b                   �m@�q�q�?             8@       \       _                    �?X�Cc�?
             ,@       ]       ^                   �l@�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        `       a                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        e       �       	          ��� @���y4F�?-             S@       f              	          033�?��h!��?#            �L@       g       ~                    �?d}h���?             E@       h       m                    �?��R[s�?            �A@        i       j                   �n@      �?             $@        ������������������������       �                     @        k       l                   �c@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        n       o                   �`@�J�4�?             9@        ������������������������       �                     �?        p       s                    �?      �?             8@        q       r                   �p@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        t       y                    �?�KM�]�?             3@       u       x       	             �?@4և���?	             ,@        v       w                   j@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        z       }       
             �?z�G�z�?             @        {       |       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@��S���?             .@       �       �                   `b@      �?              @       �       �                   p`@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             3@        �       �       
             �?�8��8��?J             ^@       �       �                    `@ ��WV�??             Z@        �       �                   @_@���y4F�?             3@       �       �                   �b@�t����?             1@       �       �                    �Q@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        0            @U@        �       �                    �?      �?             0@        �       �       	             @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   `@�B-]��?�            �q@        �       �       
             �?b1<+�C�?,            @R@       �       �                   �r@ i���t�?            �H@       �       �                   �j@���.�6�?             G@       �       �                    \@�S����?             3@        �       �                    @L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @P@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        ������������������������       �                     ;@        �       �       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    @ �q�q�?             8@       ������������������������       �                     6@        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          ����?��5���?�            �j@       �       �       
             �?L�[2[
�?{            �f@        �       �                   �b@"Ae���?            �G@        �       �                    �?�G�z��?             4@        �       �                    �?և���X�?             @        �       �                   pn@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    `P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     G@�n_Y�K�?	             *@        ������������������������       �                      @        �       �                    �?���!pc�?             &@       ������������������������       �                     @        �       �                    �?      �?             @       �       �                    ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �[@�+$�jP�?             ;@        ������������������������       �                     �?        �       �                   �d@8�Z$���?             :@        �       �       	          hff�?�	j*D�?             *@        �       �                   �o@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    c@@A��q�?_            �`@       �       �                   �^@�]���?S            �\@        ������������������������       �        %            �H@        �       �       	            �?Pa�	�?.            �P@       �       �                    �L@ �.�?Ƞ?(             N@       ������������������������       �                    �G@        �       �                    @M@$�q-�?
             *@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �       	          pff�?      �?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   Pc@ףp=
�?             4@        ������������������������       �                      @        ������������������������       �                     2@        �       �                   Ph@     ��?             @@        �       �                    d@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �e@�q�q�?             8@       �       �                    �?���N8�?             5@       �       �                    �?r�q��?             2@       ������������������������       �                     $@        �       �                    �O@      �?              @       �       �                    �?����X�?             @       ������������������������       �                     @        �       �                     H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �k@�q�q�?             @        ������������������������       �                     �?        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �B`�P4�?��ϊ�e�?`��c.�?�Ug�{�?~)]����?AkQ���?�pR���?�c+����?�lٲe˶?iҤI�&�?              �?�q�q�?�q�q�?      �?        Lg1��t�?�YLg1�?333333�?ffffff�?              �?      �?        �;�;�?��؉���?�{a���?a����?d!Y�B�?ӛ���7�?      �?      �?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?{�G�z�?���Q��?(�����?�5��P�?      �?        �$I�$I�?�m۶m��?              �?      �?      �?d!Y�B�?ӛ���7�?              �?�a�a�?=��<���?              �?�q�q�?�q�q�?      �?        �?�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?�1�c��?�s�9��?      �?              �?      �?      �?        �?�������?              �?�������?�������?              �?      �?        �������?""""""�?S�n0�?�Y7�"��?�$I�$I�?۶m۶m�?              �?      �?        ���@���?��~5&�?�������?333333�?�$I�$I�?۶m۶m�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?m�w6�;�?L� &W�?�ڕ�]��?ە�]���?<<<<<<�?�?n۶m۶�?�$I�$I�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?%I�$I��?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?              �?              �?        (������?6��P^C�?p�}��?Hp�}�?۶m۶m�?I�$I�$�?PuPu�?X|�W|��?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?        {�G�z�?�z�G��?      �?              �?      �?�������?�������?      �?                      �?(�����?�k(���?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?�������?�������?      �?      �?      �?                      �?              �?              �?�������?�?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?UUUUUU�?UUUUUU�?;�;��?O��N���?(������?6��P^C�?�?<<<<<<�?      �?      �?              �?      �?              �?              �?                      �?      �?      �?۶m۶m�?�$I�$I�?      �?                      �?              �?�d���?i6�����?Ĉ#F��?�;w�ܹ�?����X�?/�����?Y�B��?���7���?^Cy�5�?(������?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?      �?              �?      �?      �?                      �?l9��/��?Q�@��?��{��{�?�!�!�?�w6�;�?W�+���?�������?�������?�$I�$I�?۶m۶m�?333333�?�������?              �?      �?              �?      �?              �?      �?        ى�؉��?;�;��?      �?        t�E]t�?F]t�E�?              �?      �?      �?      �?      �?      �?                      �?      �?        /�����?B{	�%��?              �?;�;��?;�;��?vb'vb'�?;�;��?      �?      �?      �?      �?      �?                      �?              �?�q�q�?�q�q�?      �?                      �?      �?        ��)F�?t��:W�?��ʇq�?���ϑ?      �?        |���?|���?wwwwww�?�?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?UUUUUU�?      �?              �?      �?      �?      �?              �?      �?              �?        �������?�������?              �?      �?              �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?�a�a�?��y��y�?�������?UUUUUU�?      �?              �?      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��(.hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK酔h��B@:         v                    �?({E�B��?�           ��@              5       	          ����?T����?�            y@               4                    f@N�N����?\            @b@                                 �e@��c:�?X            @a@                                   `@`�H�/��?!            �I@                                   �L@�d�����?             3@                     
             �?�n_Y�K�?             *@       ������������������������       �                     @        	              	          @33�?����X�?             @       
                           �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @@               +       	          833�?|�|k6��?7            �U@              $                   �`@�'�=z��?*            �P@                                  �?~|z����?             �J@                     
             �?���Q��?             D@        ������������������������       �                     *@                                  e@�����H�?             ;@                                  �L@$�q-�?             :@                                  �I@ �q�q�?             8@       ������������������������       �                     0@                                  �[@      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                  `l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                !                    �?$�q-�?             *@       ������������������������       �                     &@        "       #                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       (                   �a@�	j*D�?
             *@       &       '                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        )       *                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ,       -       	          ����?؇���X�?             5@       ������������������������       �        	             (@        .       /                    �?�q�q�?             "@        ������������������������       �                      @        0       3       
             �?؇���X�?             @       1       2                   @_@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        6       E                   �\@��O���?�            �o@        7       D                    �P@������?             >@       8       C                    �L@�+$�jP�?             ;@       9       :                    �?�t����?             1@        ������������������������       �                      @        ;       <                   @Z@z�G�z�?
             .@        ������������������������       �                     @        =       >                   `_@���!pc�?             &@        ������������������������       �                     @        ?       B       	          033@և���X�?             @        @       A                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        F       G                   �Q@4�f����?�             l@        ������������������������       �                      @        H       q                   �c@���" �?�            �k@       I       b                    �?�Wv���?�             k@       J       a       	          ���@�g�y��?e            `c@       K       `       	             @���7�?H            �[@       L       ]                    c@������?G             [@       M       N                    �?���J��?B            �Y@        ������������������������       �                     8@        O       P                    �? ���J��?2            �S@        ������������������������       �                     $@        Q       R       	          033�?г�wY;�?+             Q@        ������������������������       �                     4@        S       T                   �b@ �q�q�?             H@       ������������������������       �                     =@        U       Z                   �_@�KM�]�?             3@       V       W                   `c@�IєX�?	             1@        ������������������������       �                     @        X       Y                    �P@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        [       \                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ^       _                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �F@        c       f                   �_@\#r��?             �N@        d       e                   �p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        g       p                    �?�}�+r��?            �L@       h       k                   �`@ȵHPS!�?             :@        i       j                    @L@      �?              @       ������������������������       �                     @        ������������������������       �                      @        l       m       
             �?�X�<ݺ?
             2@       ������������������������       �                     .@        n       o                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ?@        r       u                     M@և���X�?             @       s       t       	          pff�?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        w       �                    �?Ɨ�v2U�?�            �t@       x       y                    X@v��؈�?�            Pq@        ������������������������       �                     @        z       �                    �?֙S}o�?�            �p@       {       �                    @B@��n�'��?�            �m@        |       �                    @������?             A@       }       ~                    b@r�q��?             >@        ������������������������       �                     @               �                    �? ��WV�?             :@        ������������������������       �                     @        �       �                   @^@�}�+r��?             3@        �       �       	              @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   0d@lE�x�?�            �i@        �       �       
             �?X�Cc�?	             ,@        �       �                   @^@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �]@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?XNbǃ%�?z            �g@        �       �                   @a@�<ݚ�?             B@       �       �                    �?�LQ�1	�?             7@        ������������������������       �                     ,@        �       �                   �b@�q�q�?             "@        ������������������������       �                     @        �       �       
             �?      �?             @        ������������������������       �                      @        �       �                    @H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   hr@�n_Y�K�?	             *@       �       �                   pc@���!pc�?             &@       �       �                   n@�����H�?             "@        ������������������������       �                     @        �       �       	          `ff�?z�G�z�?             @        ������������������������       �                     @        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �? ���l��?a            `c@        ������������������������       �        +            �P@        �       �       	          ���@ p�/��?6            @V@       �       �                     L@�d���?5            �U@       ������������������������       �        -            �S@        �       �                    d@�<ݚ�?             "@       �       �                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ���ٿ      �?             @@        ������������������������       �                     @        �       �       	          ���@П[;U��?             =@       �       �                    @L@      �?             8@        �       �                     I@ףp=
�?	             $@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?և���X�?             ,@       �       �                   Pc@X�<ݚ�?             "@       �       �       	          ����?և���X�?             @       �       �                    �?�q�q�?             @       �       �                   r@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?z�G�z�?             @        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��X��?#             L@       �       �                   �`@��H�}�?             I@       �       �       
             �?ȵHPS!�?             :@       �       �       	          ����?HP�s��?             9@       �       �                     P@؇���X�?	             ,@       �       �                    �?$�q-�?             *@        ������������������������       �                     @        �       �                     N@ףp=
�?             $@        �       �                    ^@�q�q�?             @        ������������������������       �                     �?        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �d@      �?             8@       �       �                   �f@����X�?             5@       �       �       
             �?���y4F�?             3@       �       �                    @M@�q�q�?             (@       �       �                    �J@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B�  Ac�Zb�?`yΨ�N�?J���h�?|��O���?�Ǐ?~�?8p���?�7��Mo�?-d!Y��?�?�������?y�5���?Cy�5��?ى�؉��?;�;��?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?              �?      �?                      �?              �?              �?�2)^ �?;���C��?|��|�?|���?��sHM0�?�	�[���?333333�?�������?              �?�q�q�?�q�q�?�؉�؉�?;�;��?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?              �?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?vb'vb'�?;�;��?      �?      �?              �?      �?        �������?333333�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        �?�������?�?wwwwww�?B{	�%��?/�����?�������?�������?      �?        �������?�������?              �?t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?              �?      �?        ߼�xV4�?d��0u��?      �?        ��p"^�?��;���?/�����?�%���^�?�B!��?��{���?F]t�E�?�.�袋�?�q�q�?�q�q�?�?______�?              �?�A�A�?��-��-�?              �?�?�?              �?UUUUUU�?�������?              �?(�����?�k(���?�?�?              �?F]t�E�?]t�E�?              �?      �?              �?      �?      �?                      �?UUUUUU�?�������?      �?                      �?      �?                      �?XG��).�?��:��?      �?      �?      �?                      �?(�����?�5��P�?�؉�؉�?��N��N�?      �?      �?              �?      �?        �q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?O}Q����?b]#V�?�f����?�e����?              �?Ŀ{��(�?� 2�]�?��Ϣ��?P���:Ǻ?xxxxxx�?�?�������?UUUUUU�?              �?O��N���?;�;��?      �?        �5��P�?(�����?]t�E�?F]t�E�?      �?                      �?      �?              �?      �?              �?      �?        Y��թX�?;�S�:�?%I�$I��?�m۶m��?�������?333333�?      �?                      �?9��8���?�q�q�?              �?      �?        �uX�Q��?kP<�q�?9��8���?�q�q�?��Moz��?Y�B��?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?      �?      �?                      �?;�;��?ى�؉��?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?        �������?�������?      �?              �?      �?              �?      �?                      �?              �?-��,�?mЦm�?      �?        �G?�я�?p�\��?�:���C�?Ȥx�L��?      �?        9��8���?�q�q�?      �?      �?              �?      �?                      �?              �?      �?      �?              �?�{a���?��=���?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?r�q��?�q�q�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?              �?        �������?�������?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?%I�$I��?n۶m۶�?
ףp=
�?{�G�z�?�؉�؉�?��N��N�?{�G�z�?q=
ףp�?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?                      �?      �?              �?      �?�m۶m��?�$I�$I�?6��P^C�?(������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJx�+hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@0         �       
             �?znt��s�?�           ��@              e                   �c@H�v  w�?           {@                                 `Q@     |�?�             x@        ������������������������       �                     @               @                    �? ��P0�?�            �w@              ;                    �?4_�����?�            �q@                                  �?�����H�?}            �i@                                   @G@�d�����?             C@        	       
                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @                                   @L@r�q��?             >@        ������������������������       �                     (@                      	          033�?�E��ӭ�?             2@                                 �`@�n_Y�K�?             *@                                  �?      �?              @                                  �?      �?             @                                 �]@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               6                   hr@$�q-�?g             e@                                  @J@8~�Q��?[             c@        ������������������������       �                     A@               5                   pb@_k,D	�?H            �]@              *       	          ����?io8�?F             ]@                                  �i@      �?             D@       ������������������������       �                     >@                !                    �?      �?             $@        ������������������������       �                     �?        "       #                    �?X�<ݚ�?             "@        ������������������������       �                     �?        $       )                   �`@      �?              @       %       (                   �[@���Q��?             @       &       '                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        +       4                   @^@P�Lt�<�?.             S@       ,       1                   �]@���N8�?             E@       -       .                    �?�(\����?             D@       ������������������������       �                     >@        /       0       	             @ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        2       3                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        ������������������������       �                      @        7       :                   s@������?             1@        8       9                   �_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             (@        <       =                    �R@P�Lt�<�?4             S@       ������������������������       �        2            @R@        >       ?                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        A       J                   0`@��O5���??            �X@       B       G                    �?$�q-�?!             J@        C       F                   �d@      �?             @       D       E                     N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        H       I                   �s@��<b�ƥ?             G@       ������������������������       �                    �F@        ������������������������       �                     �?        K       P                   �h@��c:�?             G@        L       O                   @e@���y4F�?
             3@       M       N                    �?r�q��?	             2@        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     �?        Q       X                    @K@X�<ݚ�?             ;@        R       S                    �B@"pc�
�?             &@        ������������������������       �                     �?        T       W                    �F@ףp=
�?             $@        U       V                   �o@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        Y       ^       	          `ff�?      �?             0@        Z       [                    �?�����H�?             "@       ������������������������       �                     @        \       ]                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        _       `                   0b@����X�?             @        ������������������������       �                     @        a       b                   �`@      �?             @        ������������������������       �                     �?        c       d                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        f       o                    �?`�(c�?            �H@        g       j                     M@p�ݯ��?
             3@       h       i                   �r@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        k       n                   �c@����X�?             @       l       m                   @]@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        p       �       	          `ff@�������?             >@       q       r                    �A@�>4և��?             <@        ������������������������       �                     �?        s       z       	          ����?PN��T'�?             ;@        t       u                   �j@և���X�?             @        ������������������������       �                      @        v       y                   pe@���Q��?             @       w       x                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        {       �                   e@P���Q�?             4@        |       }                   Pl@      �?              @       ������������������������       �                     @        ~                          �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        �       �                    c@RB)��.�?�            �r@        �       �       	          ����?tk~X��?             B@        �       �                    �?      �?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?$�q-�?             :@       �       �                    �O@�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?        �       �                    �?      �?              @        �       �                   �[@�q�q�?             @        ������������������������       �                     �?        �       �                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��%p���?�            �p@       �       �                    \@�kb97�?�            �l@        �       �                    �?8�Z$���?            �C@        �       �                    �L@      �?             0@       �       �                   �[@�q�q�?
             .@       �       �                    �?z�G�z�?             $@        �       �                   g@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    �?      �?}             h@        �       �       	          833�?$�q-�?            �C@       ������������������������       �                    �@@        �       �                   �`@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                     L@���J��?d             c@       ������������������������       �        Q            �^@        �       �                   �c@ףp=
�?             >@       ������������������������       �                     8@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �j@ҳ�wY;�?             A@        �       �                   �d@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        �       �                    �?b�2�tk�?             2@       �       �                    @K@��
ц��?             *@       �       �                   �`@      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @       �       �                    b@z�G�z�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  ����?��}t��?�����?�_���?      �?     ��?      �?        �@ �?�~�����?ӵ8f��?FI�8S,�?�q�q�?�q�q�?y�5���?Cy�5��?      �?      �?      �?                      �?UUUUUU�?�������?              �?r�q��?�q�q�?ى�؉��?;�;��?      �?      �?      �?      �?      �?      �?              �?      �?              �?              �?                      �?              �?;�;��?�؉�؉�?�5��P�?������?              �?��c+���?����/��?GX�i��?|a���?      �?      �?              �?      �?      �?              �?r�q��?�q�q�?              �?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        (�����?���k(�?�a�a�?��y��y�?�������?333333�?              �?�������?�������?              �?      �?              �?      �?              �?      �?                      �?      �?        �?xxxxxx�?�������?�������?              �?      �?                      �?(�����?���k(�?              �?UUUUUU�?UUUUUU�?              �?      �?        ��S�r
�?�Cc}�?;�;��?�؉�؉�?      �?      �?      �?      �?              �?      �?                      �?d!Y�B�?��7��M�?              �?      �?        �7��Mo�?-d!Y��?(������?6��P^C�?UUUUUU�?�������?      �?                      �?      �?        r�q��?�q�q�?/�袋.�?F]t�E�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�q�q�?�q�q�?              �?      �?      �?              �?      �?        �m۶m��?�$I�$I�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?������?4և����?Cy�5��?^Cy�5�?UUUUUU�?�������?              �?      �?        �m۶m��?�$I�$I�?�������?UUUUUU�?              �?      �?                      �?�������?�������?�$I�$I�?�m۶m��?              �?&���^B�?h/�����?�$I�$I�?۶m۶m�?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?ffffff�?�������?      �?      �?      �?              �?      �?              �?      �?              �?                      �?S֔5eM�?���)k��?9��8���?r�q��?      �?      �?      �?                      �?;�;��?�؉�؉�?�q�q�?��8��8�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?$�q���?q��;2l�?�Y�	qV�?�cj`?;�;��?;�;��?      �?      �?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?333333�?      �?                      �?              �?      �?              �?      �?�؉�؉�?;�;��?      �?              �?      �?              �?      �?        ______�?�?      �?        �������?�������?      �?              �?      �?      �?              �?      �?              �?      �?        �������?�������?      �?      �?              �?      �?        �8��8��?9��8���?�؉�؉�?�;�;�?      �?      �?              �?۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?      �?              �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJH�SshG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKɅ�h��B@2         ~       
             �?6������?�           ��@                                 f@ęI0�?           pz@                                   �?P���Q�?P             ^@                                   �?r�q��?             (@              
                    �?�C��2(�?             &@                                  �[@      �?             @        ������������������������       �                      @               	                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   �? 7���B�?I             [@                                   ]@�r����?             .@                      	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@                                  �_@����D��?A            @W@                                   �K@ >�֕�?            �A@        ������������������������       �                     2@                                   �?�t����?             1@                                  �L@@4և���?             ,@                      	             �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             (@                                  �^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        '             M@                S                    �?l��wC�?�            �r@        !       F       	          ����?�;_��?K            @\@       "       E                   �e@��]�T��?8            �T@       #       ,                    �?��Q��?7             T@        $       %                   @_@�>����?             ;@        ������������������������       �                     $@        &       '                   �\@�t����?             1@        ������������������������       �                     �?        (       )                   pe@      �?
             0@       ������������������������       �                     ,@        *       +                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        -       .                   �_@�F�j��?&            �J@        ������������������������       �                      @        /       6       	          ����?���Q��?            �F@        0       3                   �`@8�Z$���?
             *@        1       2                   �h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        4       5                    �K@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        7       <                    �K@     ��?             @@        8       9                   �p@��S�ۿ?	             .@       ������������������������       �                     (@        :       ;                   �q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        =       >                   Pb@ҳ�wY;�?             1@        ������������������������       �                     @        ?       B                   �l@���Q��?             $@        @       A                    `P@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        C       D                     P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        G       L                   �a@�4�����?             ?@       H       K                    �?r�q��?             2@        I       J       
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        M       R                   (u@��
ц��?             *@       N       O       
             �?���|���?             &@        ������������������������       �                      @        P       Q       	             @X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        T       a                    �?�˹�m��?}            �g@        U       `                   �b@�q�q�?             8@       V       _       	          ����?���!pc�?             6@       W       \                    �?��
ц��?	             *@       X       Y                   �s@����X�?             @       ������������������������       �                     @        Z       [                     K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ]       ^                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        b       s                    �?x�}���?j            �d@       c       d                   �Z@P����?\            `b@        ������������������������       �                     �?        e       r                    �? ��֛�?[            @b@       f       o                   �b@P�Lt�<�?E            �\@       g       n                    `@ �Jj�G�?C            �[@        h       m       	          `ff�?�7��?            �C@        i       l                    �O@z�G�z�?             $@       j       k       	             �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     =@        ������������������������       �        +            �Q@        p       q                    �J@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @@        t       w                   �j@�S����?             3@        u       v                   �i@      �?             @        ������������������������       �                      @        ������������������������       �                      @        x       y                   �a@��S�ۿ?
             .@       ������������������������       �                     $@        z       {                    �?z�G�z�?             @        ������������������������       �                     @        |       }                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               �                    �K@Σq���?�            ps@       �       �                   �S@X��*"�?�            `k@        �       �                   �\@     ��?
             0@        �       �       	          @33�?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �?@���p��?�            `i@        �       �                   0j@     ��?             H@        �       �                   @c@�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   Pb@���H��?             E@       ������������������������       �                     8@        �       �                    @K@�E��ӭ�?             2@       �       �                    �?�r����?
             .@        ������������������������       �                     @        �       �                    �G@"pc�
�?             &@        ������������������������       �                     @        �       �                   �`@���Q��?             @        ������������������������       �                     �?        �       �                   �q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        d            `c@        �       �                    �?�+Fi��?:             W@       �       �                   @E@��0u���?&             N@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �N@���B���?!             J@       �       �                    �?     ��?             @@       �       �                   @Y@������?             ;@        ������������������������       �                     �?        �       �                    @N@�θ�?             :@       �       �       	          hff @؇���X�?             5@       �       �                    �?ףp=
�?             4@       �       �                    �M@r�q��?             (@       �       �                   �_@�C��2(�?             &@        �       �                   �l@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          033@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        �       �                   Pp@      �?             @@       �       �                    �?r�q��?             2@       �       �                   @b@�q�q�?             "@       �       �                   �`@؇���X�?             @        �       �       	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?X�Cc�?             ,@        �       �                   �^@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��X�5�?��S�$e�?�k���?e����?�������?ffffff�?UUUUUU�?�������?F]t�E�?]t�E�?      �?      �?              �?      �?      �?      �?                      �?              �?      �?        h/�����?	�%����?�?�������?      �?      �?              �?      �?                      �?X`��?P?���O�?�A�A�?��+��+�?              �?�?<<<<<<�?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?מ�;�C�?��b4��?��Ź��?�(�u���?KԮD�J�?jW�v%j�?�������?ffffff�?�Kh/��?h/�����?      �?        <<<<<<�?�?              �?      �?      �?      �?              �?      �?              �?      �?        ��sHM�?:�&oe�?              �?333333�?�������?;�;��?;�;��?      �?      �?              �?      �?        F]t�E�?]t�E�?              �?      �?              �?      �?�������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?        �������?333333�?333333�?�������?      �?                      �?�������?�������?              �?      �?                      �?��RJ)��?���Zk��?UUUUUU�?�������?      �?      �?      �?                      �?              �?�;�;�?�؉�؉�?]t�E]�?F]t�E�?      �?        r�q��?�q�q�?      �?                      �?              �?^Cy�5�?��P^Cy�?UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?�؉�؉�?�;�;�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        4u~�!��?�(፦�?���+ݛ?�_��!�?      �?        �P�B�
�?{��իW�?(�����?���k(�?��)A��?k߰�k�?�A�A�?��[��[�?�������?�������?�q�q�?�q�q�?              �?      �?              �?                      �?              �?      �?      �?              �?      �?                      �?^Cy�5�?(������?      �?      �?              �?      �?        �?�������?              �?�������?�������?              �?      �?      �?      �?                      �?!�J���?|_��oH�?��C2��?x��m���?      �?      �?333333�?�������?      �?                      �?              �?�W�Δ�?xÏ���?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�0�0�?��y��y�?      �?        �q�q�?r�q��?�������?�?      �?        /�袋.�?F]t�E�?      �?        333333�?�������?              �?      �?      �?      �?                      �?              �?      �?        ���,d!�?����7��?�������?""""""�?      �?      �?      �?                      �?��؉���?ى�؉��?      �?      �?B{	�%��?{	�%���?              �?ى�؉��?�؉�؉�?۶m۶m�?�$I�$I�?�������?�������?�������?UUUUUU�?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?                      �?      �?                      �?�������?333333�?      �?                      �?333333�?�������?              �?      �?        ffffff�?�������?      �?                      �?      �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?%I�$I��?�m۶m��?UUUUUU�?�������?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�8�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKӅ�h��B�4         ~       
             �?�+	G�?�           ��@              C                    �?z�G�z�?           �{@                     	          ����?�ma�H��?�             s@               	                   @l@��{H�?3            �U@                                  �?�.ߴ#�?$            �N@                                   @N@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        !             L@        
                           �?
j*D>�?             :@                                   �?      �?              @        ������������������������       �                     @                                  �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   \@�E��ӭ�?
             2@        ������������������������       �                     @                      	             �?�r����?	             .@       ������������������������       �                     "@                                  pd@�q�q�?             @                                  �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               &                    @G@F��}��?�            `k@               %                    �?6YE�t�?            �@@                                  @D@��a�n`�?             ?@        ������������������������       �                     2@                                  �Z@�θ�?	             *@        ������������������������       �                     �?               "                   �e@r�q��?             (@                !                    ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        #       $                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        '       @                   {@(��m,��?w            @g@       (       =                    �R@hl �&�?u             g@       )       <                    �?�&���?s            �f@       *       -                   `Q@`�c�г?S             _@        +       ,       
             �?r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        .       5       	          ����?������?J             \@        /       4                   Xw@���7�?             F@       0       3                   �[@ qP��B�?            �E@        1       2                   `_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     D@        ������������������������       �                     �?        6       ;                    �J@ ��ʻ��?-             Q@        7       :                   �_@@4և���?
             ,@        8       9                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �        #             K@        ������������������������       �                     �L@        >       ?                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        A       B                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        D       O                   �Q@��2�,�?Y            �`@        E       N                   �c@      �?             @@       F       G                   �c@��S�ۿ?             >@       ������������������������       �                     7@        H       M                    �?����X�?             @       I       J                     M@      �?             @        ������������������������       �                     �?        K       L       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        P       }                    �?�7i���?D            �Y@       Q       Z                    �?:�1�(��?:            @U@        R       Y                   �b@��2(&�?             6@       S       T                   p@�����?             5@       ������������������������       �        
             ,@        U       X       	             �?����X�?             @       V       W                   �c@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        [       |                   �r@X�<ݚ�?*            �O@       \       ]       
             �?>n�T��?'             M@        ������������������������       �                     @        ^       s                   a@�\�u��?#            �I@       _       j                   �l@     ��?             @@        `       a                   �e@r�q��?             (@        ������������������������       �                     �?        b       i                    �?�C��2(�?             &@       c       h                   @_@�����H�?             "@       d       e                   �[@z�G�z�?             @        ������������������������       �                      @        f       g                   �k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        k       l                   0b@      �?             4@        ������������������������       �                     @        m       r                    �?X�Cc�?             ,@       n       o                   0c@      �?              @        ������������������������       �                     @        p       q                    �E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        t       u                    @�}�+r��?             3@       ������������������������       �        	             &@        v       {                   �o@      �?              @        w       x       	          @33�?�q�q�?             @        ������������������������       �                     �?        y       z                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             1@               �       	          ����?�+�ԗ�?�            `r@       �       �                    �?�8��8��?�            �i@        �       �                    �?r٣����?            �@@        �       �                    �?�q�q�?	             (@        �       �                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    ]@      �?              @        ������������������������       �                     @        �       �                   �`@z�G�z�?             @        �       �                    _@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     L@؇���X�?             5@       ������������������������       �                     ,@        �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                   �a@      �?             @        ������������������������       �                     �?        �       �                   �m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�}�+r��?o            `e@        �       �                    �H@*
;&���?             G@       ������������������������       �                     ;@        �       �                   Pd@p�ݯ��?             3@       �       �                    �?      �?             ,@       �       �                   �g@�z�G��?             $@        ������������������������       �                     @        �       �                    �?      �?             @       �       �                    @J@���Q��?             @        ������������������������       �                      @        �       �                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �t@@�n�1�?Q            @_@       ������������������������       �        N            @^@        �       �                    �N@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?f.i��n�?;            �V@       �       �                   �c@�����?+             Q@        �       �                    `@      �?             (@        ������������������������       �                     @        �       �                    c@���Q��?             @        ������������������������       �                      @        �       �                    �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    Z@@4և���?#             L@        ������������������������       �                     �?        �       �                    @G@�1�`jg�?"            �K@        �       �                    �?z�G�z�?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          pff�?`2U0*��?             I@        �       �                   �a@      �?             0@       ������������������������       �                     (@        �       �                   �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     A@        �       �                   hp@�X����?             6@       �       �       	          `ff�?���y4F�?             3@       �       �                    @M@�8��8��?	             (@       ������������������������       �                      @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?և���X�?             @       �       �                    �?z�G�z�?             @        �       �                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  ��C�l�?z?+^���?ffffff�?ffffff�?k�k��?��G��G�?/�I���?���C���?XG��).�?�K�`m�?333333�?�������?      �?                      �?              �?;�;��?b'vb'v�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?r�q��?�q�q�?      �?        �?�������?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?����?��Ǐ?�?e�M6�d�?'�l��&�?�c�1Ƹ?�s�9��?              �?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?      �?      �?              �?      �?        �������?�������?      �?                      �?      �?        EM4�D�?�.����?Y�B��?ozӛ���?4O��I�?��ҟ��?��RJ)��?��Zk���?UUUUUU�?�������?      �?                      �?۶m۶m�?I�$I�$�?F]t�E�?�.�袋�?�}A_З?��}A�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �?�������?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?&���[�?�~5&��?      �?      �?�?�������?              �?�$I�$I�?�m۶m��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        }}}}}}�?AAAAAA�?�������?�������?��.���?t�E]t�?=��<���?�a�a�?      �?        �m۶m��?�$I�$I�?      �?      �?              �?      �?              �?                      �?�q�q�?r�q��?��{a�?,�4�rO�?      �?        �?�������?      �?      �?�������?UUUUUU�?              �?]t�E�?F]t�E�?�q�q�?�q�q�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?      �?              �?�m۶m��?%I�$I��?      �?      �?      �?              �?      �?      �?                      �?              �?(�����?�5��P�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?                      �?���X�?������?UUUUUU�?UUUUUU�?>���>�?|���?�������?�������?      �?      �?      �?                      �?      �?      �?              �?�������?�������?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �5��P�?(�����?���,d!�?8��Moz�?      �?        ^Cy�5�?Cy�5��?      �?      �?ffffff�?333333�?      �?              �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �rh��|�?����Mb�?      �?              �?      �?      �?                      �?�`�`�?�>�>��?�������?xxxxxx�?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        n۶m۶�?�$I�$I�?              �?A��)A�?�־a�?�������?�������?      �?      �?              �?      �?              �?        ���Q��?{�G�z�?      �?      �?      �?              �?      �?              �?      �?              �?        ]t�E]�?�E]t��?(������?6��P^C�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJUehG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKՅ�h��B@5         ~       
             �?
���P��?�           ��@              #                    �?P���8U�?           0z@                                   �?��+��?1            �R@                                 �a@�q�q�?             E@              
                    �?      �?             8@               	       	             �?"pc�
�?             &@                                  �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?                      	             �?�θ�?	             *@                                   �D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@                      	          ����?�����H�?             2@                                    M@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             *@                                  �Q@      �?             @@        ������������������������       �                     �?               "                    c@��a�n`�?             ?@                                 �Z@؇���X�?             <@                                   @      �?             @       ������������������������       �                     @        ������������������������       �                     �?               !                    �? �q�q�?             8@                                 �e@�nkK�?             7@       ������������������������       �                     4@                                   �g@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        $       S                    �?�LQ�1	�?�            �u@       %       (                   @R@g5���?�            �o@        &       '                    @K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        )       R                   �e@�&/�E�?�             o@       *       +                   i@�}�+r��?�            �n@        ������������������������       �        @            @[@        ,       3                   �[@��g=��?b            @a@        -       2                    �K@      �?              @       .       /                   �`@r�q��?             @        ������������������������       �                     @        0       1                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        4       5                    @J@$�q-�?[            @`@        ������������������������       �                    �E@        6       ;       	          ����?�:���??            �U@        7       :                    �?      �?              @       8       9                   �Y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        <       C                   p@l{��b��?8            �S@       =       B                    Y@`���i��?             F@        >       ?                     L@z�G�z�?             @        ������������������������       �                      @        @       A                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �C@        D       I                   �_@؇���X�?            �A@        E       F                   �^@      �?              @       ������������������������       �                     @        G       H                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        J       O                    c@�����H�?             ;@       K       L                   Ps@�nkK�?             7@       ������������������������       �                     2@        M       N                   ps@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       Q                   �c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        T       a                   0`@VP��g��?A             W@        U       `                    �?X�EQ]N�?            �E@       V       [                    �?д>��C�?             =@        W       X                   �W@�q�q�?             @        ������������������������       �                     �?        Y       Z                    \@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        \       _                    \@�nkK�?             7@        ]       ^                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �        
             ,@        b       y       	          ��� @Tt�ó��?#            �H@       c       p                   �`@X�<ݚ�?             B@       d       e                    @H@��+7��?             7@        ������������������������       �                     "@        f       m                   �b@և���X�?
             ,@       g       l                   �b@����X�?             @       h       i                     I@      �?             @        ������������������������       �                     �?        j       k                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        n       o                   `]@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        q       r                     N@�θ�?             *@        ������������������������       �                     @        s       t       	          ����?      �?             @        ������������������������       �                     �?        u       v                    `P@���Q��?             @        ������������������������       �                      @        w       x       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        z       {                    @8�Z$���?             *@        ������������������������       �                     @        |       }                   �o@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               �                    �?�^qj�{�?�            �s@        �       �                    P@�Ws�x��?B            �Y@        �       �                   �]@�c�Α�?             =@        �       �       	          ����?�eP*L��?             &@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                    �N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     M@r�q��?             2@       ������������������������       �                     &@        �       �                    c@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����>�?.            �R@        �       �                   �r@b�2�tk�?             2@       �       �                   �c@��
ц��?             *@       �       �       	          `ff�?���Q��?             $@       �       �                    �?      �?              @        �       �                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@r�q��?             @        ������������������������       �                     @        �       �                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�X�C�?!             L@       �       �                   �l@,���i�?            �D@       �       �       	          hff�?�E��ӭ�?             2@       �       �                    �?�r����?             .@       �       �                    b@"pc�
�?	             &@       �       �                   Pl@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     7@        �       �                   Pe@������?             .@       �       �                   �a@8�Z$���?             *@        ������������������������       �                     @        �       �                   r@����X�?             @        �       �                   �l@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��-#���?y            �j@        �       �       	          ����? qP��B�?.            �U@       �       �                    @L@��ɉ�?!            @P@       ������������������������       �                     N@        �       �                   @d@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        �       �                    c@�? Da�?K            �_@        �       �                    �?�eP*L��?             &@        ������������������������       �                      @        �       �                   �`@�q�q�?             "@        ������������������������       �                      @        �       �                     P@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ���@t��%�?E            �\@       �       �                   �^@�g+��@�?C            �[@        ������������������������       �                    �E@        �       �                    @L@ДX��?(             Q@       ������������������������       �                    �J@        �       �                    �?��S���?
             .@       �       �                   �_@�q�q�?             (@        ������������������������       �                     @        �       �                    @M@      �?              @       �       �                   �i@z�G�z�?             @        ������������������������       �                      @        �       �                    �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �P@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�b�       h�h)h,K ��h.��R�(KK�KK��hb�BP  փmM���?>IY�8�?S(*	[�?:�u�=��?�S�n�?*�Y7�"�?UUUUUU�?UUUUUU�?      �?      �?/�袋.�?F]t�E�?�������?�������?      �?                      �?              �?�؉�؉�?ى�؉��?      �?      �?              �?      �?                      �?�q�q�?�q�q�?�������?333333�?      �?                      �?              �?      �?      �?              �?�c�1��?�s�9��?۶m۶m�?�$I�$I�?      �?      �?              �?      �?        �������?UUUUUU�?�Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?Y�B��?��Moz��?�I��6�?Ė��+��?�������?�������?              �?      �?        �s�9�?2�c�1�?(�����?�5��P�?              �?��v`��?�(�3J��?      �?      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        ;�;��?�؉�؉�?              �?��֡�l�?A&�dR�?      �?      �?�������?�������?              �?      �?                      �?�&��jq�?${�ґ�?F]t�E�?F]t�E�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?              �?      �?        �q�q�?�q�q�?d!Y�B�?�Mozӛ�?              �?�������?�������?      �?                      �?      �?      �?      �?                      �?      �?        -d!Y��?�Mozӛ�?qG�wĽ?w�qG�?|a���?a���{�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?        d!Y�B�?�Mozӛ�?      �?      �?      �?                      �?              �?              �?/�����?h�����?r�q��?�q�q�?zӛ����?Y�B��?      �?        �$I�$I�?۶m۶m�?�$I�$I�?�m۶m��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?        �؉�؉�?ى�؉��?              �?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?      �?        ���?�����?���VC�?��R�y�?�{a���?5�rO#,�?]t�E�?t�E]t�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?�������?              �?۶m۶m�?�$I�$I�?              �?      �?        �u�)�Y�?���L�?9��8���?�8��8��?�;�;�?�؉�؉�?�������?333333�?      �?      �?      �?      �?              �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?�m۶m��?%I�$I��?�����?8��18�?�q�q�?r�q��?�������?�?/�袋.�?F]t�E�?�������?�������?      �?                      �?              �?      �?                      �?      �?        wwwwww�?�?;�;��?;�;��?      �?        �m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?                      �?��sH�?�琚`��?��}A�?�}A_З??�?��? �����?      �?        333333�?�������?              �?      �?              �?        �������?AA�?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?                      �?�(�j��?�q�.�|�?���+c��?Nq��$�?      �?        �������?ZZZZZZ�?      �?        �?�������?�������?�������?              �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�)�rhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@0         j                    �?8}�ý�?�           ��@              U                    �?�����?           �{@              F       	          033�?^;|��?�            Pv@              '       
             �?�ap��?�            `t@                      	          ����?r�����?6            @V@                                   �?�����?            �H@       ������������������������       �                     =@                                  �`@      �?             4@       	       
                    �?�	j*D�?             *@        ������������������������       �                     @        ������������������������       �                     "@                                  `a@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?��Q��?             D@                                  xp@�KM�]�?             3@                                  b@r�q��?
             (@                                 p@�C��2(�?	             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?և���X�?             5@                                  `]@      �?              @        ������������������������       �                     �?                      	          ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @               "                   �l@��
ц��?             *@               !                   �c@؇���X�?             @                                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        #       &                   @`@r�q��?             @        $       %                     L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        (       =                    �? 1�/Gu�?�            �m@        )       8       	          ����?      �?#             J@       *       7       	          833�?R���Q�?             D@       +       ,                   �b@�MI8d�?            �B@        ������������������������       �                     1@        -       2                   `\@�z�G��?             4@        .       /                   �n@�q�q�?             @       ������������������������       �                     @        0       1                   �[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        3       4                    s@؇���X�?
             ,@       ������������������������       �                      @        5       6                   `s@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        9       :                    �?�q�q�?             (@        ������������������������       �                     @        ;       <       	             �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        >       ?                    @L@ S5W�?t             g@       ������������������������       �        b            `c@        @       E                   b@(;L]n�?             >@        A       D                   �_@$�q-�?             *@        B       C                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     1@        G       L                    @H@�חF�P�?             ?@        H       K                    �?���Q��?             @       I       J                   �u@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        M       P                    �?$�q-�?             :@        N       O                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        Q       R                    @���7�?             6@       ������������������������       �        
             2@        S       T                     K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        V       ]       	          033�?��X��?0             U@       W       Z       
             �?z�J��?            �G@       X       Y                    �?���}<S�?             7@        ������������������������       �                      @        ������������������������       �                     5@        [       \                   �U@�8��8��?             8@        ������������������������       �                      @        ������������������������       �                     6@        ^       i                   8r@�L���?            �B@       _       b                    �J@�X�<ݺ?             B@        `       a                   �_@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        c       d                   �c@�g�y��?             ?@       ������������������������       �                     ;@        e       f                    �N@      �?             @        ������������������������       �                      @        g       h       	          ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        k       �       
             �?�׺W4�?�            Pr@       l       �                   �b@������?�            �n@       m       �                   �e@\I���?�?�             m@       n       �                   `\@�`z����?�            `l@        o       ~       	             �?,���i�?-            �T@        p       w                   �Y@��a�n`�?             ?@       q       r                    �?�����?             5@       ������������������������       �        
             0@        s       t                    �K@���Q��?             @        ������������������������       �                      @        u       v                    �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        x       }                   �[@      �?             $@       y       z                     M@r�q��?             @        ������������������������       �                     @        {       |                   `a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               �                   �c@�IєX�?            �I@       ������������������������       �                    �C@        �       �                    �?      �?             (@       �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @����=O�?a             b@       �       �                    @L@@ݚ)�?`             b@        �       �                   �a@�"w����?/             S@       ������������������������       �        %             P@        �       �                   @Z@�8��8��?
             (@        �       �                   Pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�IєX�?1             Q@        �       �                   �q@����X�?             @       ������������������������       �                     @        �       �                   @_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�]0��<�?,            �N@       �       �                    \@�}�+r��?             C@        �       �       	             @���Q��?             @       �       �                   �^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �@@        ������������������������       �                     7@        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �H@X�Cc�?
             ,@        �       �                     D@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   `c@؇���X�?             @        �       �                   0p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��C���?            �G@        ������������������������       �                     @        �       �                    �?�q�q�?             E@       �       �                    @N@�(�Tw��?            �C@       �       �                   �c@����"�?             =@       �       �       	          033�?
j*D>�?             :@       �       �       	             �?�q�q�?             5@       �       �                   �d@��
ц��?             *@       �       �                   `m@      �?              @       �       �                    �M@�q�q�?             @       �       �                    b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  a[ӿc�?PR Np�?G-B���?q�{���?���?�����?�T�;^l�?ìF�N�?��g<��?1�9�a�?����X�?^N��)x�?              �?      �?      �?;�;��?vb'vb'�?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?�������?ffffff�?�k(���?(�����?�������?UUUUUU�?]t�E�?F]t�E�?      �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?�;�;�?�؉�؉�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?��v��?(�X�>�?      �?      �?333333�?333333�?��L���?L�Ϻ��?      �?        ffffff�?333333�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?�m۶m��?�$I�$I�?              �?      �?        <����?@bw�#v?      �?        �������?�?�؉�؉�?;�;��?      �?      �?              �?      �?              �?              �?        ��RJ)��?�Zk����?333333�?�������?      �?      �?      �?                      �?              �?;�;��?�؉�؉�?      �?      �?              �?      �?        F]t�E�?�.�袋�?              �?      �?      �?              �?      �?        %I�$I��?n۶m۶�?AL� &W�?}g���Q�?d!Y�B�?ӛ���7�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        L�Ϻ��?}���g�?�q�q�?��8��8�?�������?�������?              �?      �?        �B!��?��{���?              �?      �?      �?              �?      �?      �?              �?      �?              �?        gB����?:f���M�?������?�|����?�rO#,��?��{a�?��gG�?�s���?8��18�?�����?�s�9��?�c�1��?�a�a�?=��<���?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�?�?              �?      �?      �?      �?      �?              �?      �?                      �?��RA�/�?U��K��?r�qǡ?9��8���?(�����?Cy�5��?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�?�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?;ڼOqɠ?\2�h��?(�����?�5��P�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?      �?        333333�?�������?              �?      �?        �m۶m��?%I�$I��?�$I�$I�?۶m۶m�?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?g���Q��?L� &W�?      �?        UUUUUU�?UUUUUU�?� � �?�o��o��?�i��F�?	�=����?;�;��?b'vb'v�?UUUUUU�?UUUUUU�?�;�;�?�؉�؉�?      �?      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?      �?                      �?�������?�������?              �?      �?                      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX"4qhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@0                              �?P|�z��?�           ��@                                   �?���lv	�?l            �e@                                  �a@~h����?%             L@                     	          ����?��]�T��?            �D@              
                    �?8�Z$���?             :@              	                   �_@H%u��?             9@                                 �i@�θ�?             *@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     (@        ������������������������       �                     �?                                  0c@������?             .@       ������������������������       �        	             "@                                   �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @                      
             �?��S�ۿ?
             .@       ������������������������       �                     (@                                  �s@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �K@H��ԛ�?G            �]@       ������������������������       �        8            �W@                                  a@z�G�z�?             9@        ������������������������       �                     &@                                   �?X�Cc�?	             ,@        ������������������������       �                     @                      
             �?ףp=
�?             $@                                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        !       z       
             �?�&!��?`           x�@       "       [                    �?��E�B��?�            �t@       #       V                    �?<I����?�            �n@       $       U                   �a@�^����?n            �d@       %       H                    �?T&ss��?V            �`@       &       ?                   pb@d/
k�?D             [@       '       4                   @^@x��B�R�?;            �V@        (       +                    �?$�q-�?             :@        )       *                   `@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ,       -                    �K@���N8�?             5@        ������������������������       �                     &@        .       /       
             �?ףp=
�?             $@        ������������������������       �                      @        0       3                    �M@      �?              @        1       2                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        5       6                    �? ����?,            @P@        ������������������������       �                     1@        7       >                   �[@@��8��?!             H@        8       9                    �?�C��2(�?             &@        ������������������������       �                      @        :       ;                    @K@�����H�?             "@        ������������������������       �                     @        <       =                   �Z@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �B@        @       G                   �`@��.k���?	             1@       A       B       	          ����?      �?             (@        ������������������������       �                     @        C       D       	          ����?      �?             @        ������������������������       �                      @        E       F                    \@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        I       N       	             �?l��
I��?             ;@        J       K                   �k@�q�q�?             (@        ������������������������       �                     @        L       M                   `^@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        O       T                    `@z�G�z�?
             .@        P       S       
             �?      �?             @       Q       R                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @@        W       Z                   �`@�Fǌ��?2            �S@        X       Y                   p`@������?             B@       ������������������������       �                    �A@        ������������������������       �                     �?        ������������������������       �                    �E@        \       i                    �?rp��P��?2            �T@        ]       `                    �K@և���X�?             <@        ^       _                   �`@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        a       f                    �O@����X�?             5@       b       e                    �?@4և���?             ,@       c       d       
             �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        g       h                   �n@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        j       w                    �?"pc�
�?!            �K@        k       p       	          ����?�û��|�?             7@        l       o                   `X@r�q��?             (@        m       n                    d@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        q       r                   �[@���|���?             &@        ������������������������       �                      @        s       t       	             �?�<ݚ�?             "@       ������������������������       �                     @        u       v                   �^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        x       y                   @e@      �?             @@       ������������������������       �                     ?@        ������������������������       �                     �?        {       �                    �?�����?�            �l@       |       �       	          ����?*���?y             i@       }       �                    `R@ ��Ou��?[            �c@       ~       �                   `\@�kb97�?Z            @c@               �                    �?�>4և��?             <@       �       �                    �?���B���?             :@       �       �                    �?"pc�
�?
             6@        ������������������������       �                      @        �       �                   `l@ףp=
�?	             4@       ������������������������       �                     &@        �       �                   @Z@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    @L@�Ń��̧?L            �_@       �       �                    `@@䯦s#�?A            �Z@        �       �                    �I@��Y��]�?            �D@       ������������������������       �                     8@        �       �                    @J@�IєX�?             1@        �       �                    _@z�G�z�?             @        ������������������������       �                     @        �       �                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �        &            @P@        �       �                    �L@ףp=
�?             4@        �       �                   �a@�q�q�?             @        ������������������������       �                      @        �       �                    `@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                      @        �       �                    �?F�����?            �F@       �       �                   �c@�q�q�?             8@        ������������������������       �                     @        �       �                    b@���N8�?             5@       �       �                    @L@�n_Y�K�?	             *@       �       �                   �_@؇���X�?             @        �       �                   �g@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �p@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �`@���N8�?             5@        �       �       	          033�?؇���X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        �       �                    T@П[;U��?             =@        �       �       	             п�θ�?	             *@        ������������������������       �                      @        �       �                   0a@�C��2(�?             &@       ������������������������       �                     @        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?     ��?             0@       ������������������������       �        
             &@        �       �                   @p@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  ��erd��?;���7�?�bSi��?L�w�Z��?�m۶m��?%I�$I��?KԮD�J�?jW�v%j�?;�;��?;�;��?)\���(�?���Q��?ى�؉��?�؉�؉�?              �?      �?              �?                      �?�?wwwwww�?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        _̧^̧�?:�:��?      �?        �������?�������?      �?        %I�$I��?�m۶m��?              �?�������?�������?      �?      �?      �?                      �?      �?        S֔5eM�?֔5eMY�?AL� &W�?�l�w6��?�M!д?f�_��e�?W��1 �?ՃF��[�?= Y���?�)F�?/�����?�Kh/���?��?�����?;�;��?�؉�؉�?�������?�������?              �?      �?        �a�a�?��y��y�?              �?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �? �����? �����?              �?UUUUUU�?UUUUUU�?F]t�E�?]t�E�?              �?�q�q�?�q�q�?              �?�������?�������?              �?      �?                      �?�?�������?      �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?      �?        h/�����?Lh/����?�������?�������?              �?�m۶m��?�$I�$I�?              �?      �?        �������?�������?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?�3���?1���M��?�q�q�?�q�q�?              �?      �?                      �?�7�:���?>�b���?۶m۶m�?�$I�$I�?۶m۶m�?�$I�$I�?              �?      �?        �$I�$I�?�m۶m��?�$I�$I�?n۶m۶�?F]t�E�?]t�E�?      �?                      �?              �?�m۶m��?�$I�$I�?      �?                      �?F]t�E�?/�袋.�?��,d!�?8��Moz�?UUUUUU�?�������?�������?333333�?      �?                      �?              �?]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �@�V���?�����a�?^��C��?��s��2�?.��-���?�i�i�?�Y�	qV�?�cj`?�$I�$I�?�m۶m��?��؉���?ى�؉��?/�袋.�?F]t�E�?              �?�������?�������?      �?        9��8���?�q�q�?              �?      �?              �?      �?              �?      �?              �?        ��<��<�?�a�a�?R����?�x+�R�?8��18�?������?      �?        �?�?�������?�������?      �?              �?      �?      �?                      �?      �?              �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?؂-؂-�?�>�>��?UUUUUU�?UUUUUU�?              �?�a�a�?��y��y�?;�;��?ى�؉��?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �a�a�?��y��y�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?�{a���?��=���?�؉�؉�?ى�؉��?      �?        F]t�E�?]t�E�?              �?      �?      �?      �?                      �?      �?      �?      �?        �������?333333�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ;�3whG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKυ�h��B�3         �                    �?"�\�&U�?�           ��@              =                    �?fmCNT3�?           �y@                                  P`@��{r٣�?]            �`@                      
             �?^l��[B�?'             M@                                 �k@@-�_ .�?            �B@       ������������������������       �                     <@               
                   �`@�<ݚ�?             "@               	                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                      	          ����?�G��l��?             5@        ������������������������       �                     @                                  `X@����X�?             ,@       ������������������������       �                     $@        ������������������������       �                     @                       
             �?؀�:M�?6            �R@                                   �?l��
I��?             ;@                                  �p@r�q��?             @        ������������������������       �                     @                                  pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                    L@؇���X�?             5@       ������������������������       �        	             ,@                                   �M@և���X�?             @                                  �L@      �?             @        ������������������������       �                      @                                  p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        !       "                   `Z@��k=.��?%            �G@        ������������������������       �                     �?        #       ,                    �?�㙢�c�?$             G@        $       +                   �e@z�G�z�?
             .@       %       *                   d@      �?              @       &       )                    ^@r�q��?             @        '       (                    q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        -       6                    �?�חF�P�?             ?@       .       5                   0k@$�q-�?             :@        /       0                   �^@����X�?             @        ������������������������       �                     @        1       4       	             �?�q�q�?             @       2       3                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        7       :                    �?���Q��?             @       8       9                    ]@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ;       <       	          :33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        >       k       
             �?f��N�&�?�            �q@        ?       j                   hr@k��9�?8            �V@       @       K                    �?Ї?��f�?7            @U@        A       J       	          ����?� �	��?             9@       B       E       	          ����?b�2�tk�?             2@       C       D                    @K@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        F       I                   �l@�����H�?             "@        G       H                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        L       S                   �^@^n����?'             N@        M       R                   �b@      �?
             0@        N       O       	          ����?����X�?             @        ������������������������       �                     @        P       Q                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        T       Y                    �?�zv�X�?             F@        U       X                   �_@"pc�
�?             &@        V       W                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        Z       c                   �c@r٣����?            �@@       [       \                    �?���}<S�?             7@       ������������������������       �        
             .@        ]       b                    �?      �?              @       ^       a                    �?؇���X�?             @        _       `                   `d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        d       i                    @O@���Q��?             $@       e       f                   �]@z�G�z�?             @        ������������������������       �                      @        g       h                    c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        l       �                    @�0p<���?x             h@       m       r                    @L@x/ ��?p            �f@       n       q                   `R@�e���@�?^            @c@        o       p                    @H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        \            �b@        s       �       	          833@      �?             <@       t       u                   �^@�<ݚ�?             ;@        ������������������������       �                      @        v       �                   �d@�����?             3@       w       ~                   Hp@      �?             0@       x       }                    �?      �?	             (@       y       z                   �a@�z�G��?             $@       ������������������������       �                     @        {       |                   `c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               �                    �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �h@"pc�
�?             &@        ������������������������       �                     @        �       �                   Pl@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   Hq@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?|S��?�            �s@        �       �                    �?����e��?            �@@       �       �                   xt@������?             ;@       �       �                    �?�IєX�?             1@       ������������������������       �        	             (@        �       �                     M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    `@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pl@$�q-�?�            �q@       �       �                    �D@XB���?\             b@        �       �                    �C@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?`��(�?V            �`@       �       �                   `_@�6H�Z�?I            @]@       ������������������������       �        ,            �P@        �       �                   `]@p���?             I@        ������������������������       �                     �?        ������������������������       �                    �H@        �       �                   �]@�X�<ݺ?             2@        �       �                    @N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        �       �                   �l@L�
�$�?T            �a@        �       �                    �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   ``@DS���|�?Q             a@        �       �       	          ����?�+$�jP�?!             K@        ������������������������       �                     &@        �       �                   �^@>��C��?            �E@        �       �                   �m@ףp=
�?             4@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             (@        �       �                   `\@�LQ�1	�?             7@        ������������������������       �                     @        �       �                   `n@r�q��?             2@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    `@      �?
             0@        �       �                    @J@      �?             @        ������������������������       �                     �?        �       �                     O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?��`qM|�?0            �T@       �       �                    �Q@�:�]��?            �I@       �       �                    �?@9G��?            �H@       �       �       	          ����?����?�?            �F@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     E@        �       �       	          `ff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��j��`�?:�J;�O�?R��d��?�[��6��?�l��&��?��&�l��?��=���?�=�����?к����?S�n0E�?              �?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?1�0��?��y��y�?      �?        �$I�$I�?�m۶m��?              �?      �?        E>�S��?v�)�Y7�?h/�����?Lh/����?�������?UUUUUU�?      �?              �?      �?      �?                      �?�$I�$I�?۶m۶m�?              �?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?      �?                      �?              �?g���Q��?br1���?              �?�7��Mo�?d!Y�B�?�������?�������?      �?      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?        �Zk����?��RJ)��?�؉�؉�?;�;��?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�K�V��?ǬӢ�~�?[�[��?�'}�'}�?�������?�������?�Q����?)\���(�?9��8���?�8��8��?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        DDDDDD�?�������?      �?      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�袋.��?��.���?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        |���?>���>�?d!Y�B�?ӛ���7�?              �?      �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?        333333�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��3-�?�O�l.�?��j��j�?�Q�Q�?qV~B���?�cj`?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?9��8���?�q�q�?      �?        Q^Cy��?^Cy�5�?      �?      �?      �?      �?ffffff�?333333�?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?              �?                      �?/�袋.�?F]t�E�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        o
M`x�?�^��0}�?6�d�M6�?e�M6�d�?{	�%���?B{	�%��?�?�?              �?�������?�������?              �?      �?        333333�?�������?      �?                      �?      �?        ;�;��?�؉�؉�?�{a���?GX�i���?333333�?ffffff�?              �?      �?        t��:W�?j�����?���?�������?              �?{�G�z�?\���(\�?      �?                      �?�q�q�?��8��8�?      �?      �?      �?                      �?              �?{�e�ݾ?qJ��O$�?      �?      �?      �?                      �?�uy)�?I�ܺ�?B{	�%��?/�����?              �?qG�w��?$�;��?�������?�������?      �?      �?              �?      �?                      �?d!Y�B�?Nozӛ��?      �?        UUUUUU�?�������?      �?      �?              �?      �?              �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?��k���?�@	o4u�?�?}}}}}}�?9/���?������?l�l��?��I��I�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�3hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKӅ�h��B�4         T                   a@U�ք�?�           ��@               /       	          ����?>T���?�            �u@                                  �a@(8of��?U            `a@                                   �?8�Z$���?"             J@                     
             �?r٣����?            �@@                                  �?���N8�?             5@       ������������������������       �        
             1@                                   �?      �?             @       	       
                    \@�q�q�?             @        ������������������������       �                     �?                                   @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                   �?�q�q�?             (@                      	          433�?      �?             @       ������������������������       �                      @        ������������������������       �                      @                                   �P@      �?              @                                  \@r�q��?             @        ������������������������       �                      @                                  @Z@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@                                    @K@l�Ӑ���?3            �U@                     
             �?,���i�?            �D@                                    F@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �@@        !       $                   pk@      �?             G@        "       #       	          ����?z�G�z�?             .@       ������������������������       �                     (@        ������������������������       �                     @        %       *       	          ����?f���M�?             ?@       &       '                   @Z@�\��N��?             3@        ������������������������       �                     @        (       )       
             �?�	j*D�?             *@        ������������������������       �                     @        ������������������������       �                     "@        +       .                    ]@�8��8��?             (@        ,       -                     L@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        0       7                    �?�#-���?�            @j@        1       2       	             �?��.k���?             1@        ������������������������       �                     @        3       6                   �\@"pc�
�?             &@        4       5                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        8       O       	          pff�?�-j'�?v             h@       9       <                   �X@��a�n`�?<            @W@        :       ;                   �W@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        =       N                    �?�+Ĺ+�?6            �T@       >       K       
             �?��2(&�?             F@       ?       J                    �Q@��(\���?             D@       @       C                    �?�7��?            �C@        A       B       
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        D       E                    _@Pa�	�?            �@@       ������������������������       �                     8@        F       I                   �_@�����H�?             "@        G       H                   �_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        L       M                    �I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        P       Q                    s@ �ׁsF�?:             Y@       ������������������������       �        5            �V@        R       S                    t@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        U       �                    �?��<:J�?�            x@        V       �                   �e@Lv���?X            @a@       W       |       	          033�?�F.< �?S            �`@       X       y                    �N@=��T�?*            �Q@       Y       r       	          833�?����5�?$            �N@       Z       a       
             �?������?            �F@        [       \                    �?�nkK�?             7@       ������������������������       �        	             2@        ]       `                    @J@z�G�z�?             @       ^       _                   pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        b       q                    s@      �?             6@       c       d                   �b@D�n�3�?             3@        ������������������������       �                     @        e       p                    a@������?
             .@       f       o       	          ����?���|���?             &@       g       h                    �?X�<ݚ�?             "@        ������������������������       �                     @        i       j                    �?r�q��?             @        ������������������������       �                      @        k       l                    �?      �?             @        ������������������������       �                     �?        m       n                    @K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        s       x                    �?      �?	             0@       t       u                    X@���!pc�?             &@        ������������������������       �                      @        v       w                   q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        z       {                     R@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        }       �                   Pe@`Jj��?)             O@       ~       �                   Pa@P���Q�?'             N@               �       	          033@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �M@h�����?%             L@        �       �                    m@�����?             5@        ������������������������       �        	             &@        �       �                   @n@z�G�z�?	             $@        ������������������������       �                     �?        �       �                   r@�����H�?             "@        �       �       	             �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �A@        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �K@Ƴ���?�            �n@       �       �       
             �?�������?u             g@        �       �                   �d@���|���?            �K@       �       �                     J@�\��N��?             C@       �       �                    �?����X�?             5@        �       �                    b@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        �       �                    �?@�0�!��?	             1@        ������������������������       �                     @        �       �                    �J@�z�G��?             $@        ������������������������       �                     @        �       �                    �?      �?             @       �       �                   �c@      �?             @       �       �                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �       	          ����?�t����?             1@        ������������������������       �                     �?        �       �                   �k@      �?
             0@        ������������������������       �                     $@        �       �                   �[@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   pf@��G^�C�?V            @`@       ������������������������       �        G             Z@        �       �                   �S@ ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                    �?�P�*�?"             O@        �       �       
             �?      �?             0@        ������������������������       �                     �?        ������������������������       �                     .@        �       �                    �?(옄��?             G@        �       �                    _@�q�q�?             (@        �       �                   Pn@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �m@      �?              @        �       �                    �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     O@h+�v:�?             A@       �       �                    @�GN�z�?             6@       �       �                   �c@������?
             .@        �       �                   �a@ףp=
�?             $@        �       �                    �M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ��� @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	           33@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   n@�q�q�?             (@        ������������������������       �                     @        �       �       
             �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B0  ᓔ��?�5�;��?
�a��,�?>�'R�4�?Fΰ�R��?ݘ��V��?;�;��?;�;��?|���?>���>�?�a�a�?��y��y�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?�������?�������?      �?      �?      �?                      �?      �?      �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?�7[�~��?/�I���?�����?8��18�?      �?      �?      �?                      �?      �?              �?      �?�������?�������?              �?      �?        ��RJ)��?��Zk���?�5��P�?y�5���?              �?vb'vb'�?;�;��?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        _�_�?�A�A�?�?�������?      �?        F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?                      �?              �?�1�K��?��LF�W�?�c�1Ƹ?�s�9��?333333�?ffffff�?              �?      �?        ���ˊ��?(፦ί�?t�E]t�?��.���?333333�?�������?�A�A�?��[��[�?UUUUUU�?�������?      �?                      �?|���?|���?              �?�q�q�?�q�q�?      �?      �?      �?                      �?              �?      �?              �?      �?              �?      �?                      �?{�G�z�?�G�z��?              �?�q�q�?�q�q�?      �?                      �?E��޲�?v���C��??���(�?w`��k�?>����?|��|�?�������?�:��:��?������?��).��?�?wwwwww�?d!Y�B�?�Mozӛ�?              �?�������?�������?      �?      �?              �?      �?                      �?      �?      �?(������?l(�����?      �?        �?wwwwww�?F]t�E�?]t�E]�?�q�q�?r�q��?      �?        UUUUUU�?�������?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?              �?      �?F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?                      �?              �?9��8���?�q�q�?      �?                      �?�B!��?���{��?�������?ffffff�?      �?      �?              �?      �?        �$I�$I�?�m۶m��?�a�a�?=��<���?              �?�������?�������?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?              �?      �?      �?      �?                      �?      �?        ���2��?����4[�?��y�^�?��1�8�?]t�E]�?F]t�E�?y�5���?�5��P�?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?ZZZZZZ�?�������?      �?        ffffff�?333333�?      �?              �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?<<<<<<�?�?              �?      �?      �?      �?        �������?UUUUUU�?              �?      �?        �����? ����?      �?        O��N���?;�;��?              �?      �?        �RJ)���?�Zk����?      �?      �?              �?      �?        ӛ���7�?���,d�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        xxxxxx�?�������?]t�E�?�袋.��?�?wwwwww�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ� �NhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK݅�h��B@7         v                    �?�!���?�           ��@              E       
             �?���Jt��?�            �w@              (       	             �?�.�.���?�            Pq@                      	          833�?Ί��2�?\            �`@        ������������������������       �        %             I@               !                   �a@\`*�s�?7             U@                                   �?     ��?*             P@                                  �?r�q��?             H@        	       
                   �Z@      �?	             (@        ������������������������       �                     �?                                   �?"pc�
�?             &@                                  �c@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                  0a@*O���?             B@                                 �t@����X�?             <@                                 �e@D�n�3�?             3@        ������������������������       �                     @                                  �q@�q�q�?             (@                                  @K@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@                                   �?      �?              @                                  _@      �?             @        ������������������������       �                      @                                   �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     0@        "       '                    �?P���Q�?             4@       #       $                   @e@ףp=
�?             $@       ������������������������       �                     @        %       &                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        )       4       
             �?��LsƔ�?_            �a@        *       1                   �r@`Jj��?             ?@       +       0                    �?XB���?             =@        ,       /                   �T@      �?             @       -       .                   @^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     9@        2       3                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        5       B                    �Q@h�����?J             \@       6       =                   pb@Ц�f*�?H            �[@       7       <                   �\@�K}��?@            �Y@        8       ;                   �`@      �?             @        9       :                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        <            �X@        >       A                   �a@      �?              @        ?       @                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        C       D                   `g@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        F       U                    �?�ǧ\�?D            �Z@        G       P                     N@*;L]n�?             >@       H       O                   �b@      �?             0@       I       N                     H@؇���X�?
             ,@        J       M       	          ����?�q�q�?             @       K       L                     D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        Q       T                    �?@4և���?             ,@        R       S                   0c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        V       Y                    �?�����?2             S@        W       X                   �d@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        Z       m                    �?�y(dD�?+            @P@       [       h                   pc@���� �?            �D@       \       a       	          ����?�חF�P�?             ?@       ]       `                   @E@`2U0*��?             9@        ^       _       	          @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        b       c       	             �?�q�q�?             @        ������������������������       �                     @        d       g                    �?�q�q�?             @       e       f                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        i       j                     H@���Q��?             $@        ������������������������       �                     @        k       l                   �m@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        n       q       	          033�?      �?             8@       o       p                    h@      �?
             0@       ������������������������       �                     $@        ������������������������       �                     @        r       s                   �_@      �?              @        ������������������������       �                     �?        t       u                    �K@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        w       �                   �c@�-����?�            �u@        x       �                    �?�<ݚ�?            �F@       y       z       
             �?�n_Y�K�?             :@        ������������������������       �                     �?        {       �                   �b@���Q��?             9@       |       �                   �c@�eP*L��?             6@       }       ~       	             п�t����?             1@        ������������������������       �                     @               �                   �Q@؇���X�?
             ,@       �       �                    _@$�q-�?	             *@       �       �                    �?z�G�z�?             @        �       �                    \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@        �       �       
             �?0z���?�             s@        �       �                    �?���o� �?D            �Y@       �       �       	          033�?�i#[��?8             U@       �       �                   �l@h�����?'             L@        �       �                   �b@     ��?             0@       �       �                   �j@$�q-�?             *@       ������������������������       �                     @        �       �                   �\@؇���X�?             @        ������������������������       �                      @        �       �                   �^@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   pi@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�G�z��?             D@        �       �                    �?�	j*D�?
             *@        ������������������������       �                     @        �       �                   Po@      �?              @       �       �                   �a@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �p@�q�q�?             ;@       �       �                    �?r�q��?	             2@       �       �                   b@�<ݚ�?             "@        ������������������������       �                     @        �       �       
             �?���Q��?             @        ������������������������       �                     �?        �       �                   �c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �L@�����H�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �`@�q�q�?             "@        ������������������������       �                     @        �       �                   �r@      �?             @        ������������������������       �                      @        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �n@X�Cc�?             <@       �       �                   Pm@     ��?
             0@       �       �                   pb@���|���?	             &@       �       �                   �j@�<ݚ�?             "@        �       �                    @�q�q�?             @       �       �                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    e@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �h@�KM�]�?             3@        ������������������������       �                      @        ������������������������       �                     1@        �       �                    �? �u%���?�            `i@        �       �                    �?���7�?             6@       ������������������������       �                     (@        �       �                    �?ףp=
�?             $@        �       �                   �k@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Hp@@�:;��?o            �f@       ������������������������       �        R            �`@        �       �                    _@��<b�ƥ?             G@        �       �                   @b@�IєX�?
             1@        �       �                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     =@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  v��W�?E�q���?����Fj�?�Y�In%�?���o+ͺ?���Z��?���[��?���?              �?b�a��?��<��<�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?�q�q�?�$I�$I�?�m۶m��?(������?l(�����?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?      �?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?�������?ffffff�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?-)D�{�?m���G��?�B!��?���{��?�{a���?GX�i���?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?      �?                      �?�$I�$I�?�m۶m��?�־a�?!O	� �?�?�������?      �?      �?      �?      �?      �?                      �?              �?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?�&oe��?���!5��?�������?""""""�?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?                      �?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?Q^Cy��?^Cy�5�?]t�E�?F]t�E�?      �?                      �?�J��J��?Wj�Vj��?jW�v%j�?,Q��+�?�Zk����?��RJ)��?���Q��?{�G�z�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �������?333333�?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?        �r},(�?��ů�?�q�q�?9��8���?ى�؉��?;�;��?              �?�������?333333�?]t�E�?t�E]t�?�������?�������?      �?        �$I�$I�?۶m۶m�?;�;��?�؉�؉�?�������?�������?      �?      �?              �?      �?                      �?              �?      �?              �?                      �?              �?�.��.��?�D�D��?C���?r^�	��?��<��<�?�a�a�?n۶m۶�?%I�$I��?      �?      �?�؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?vb'vb'�?;�;��?      �?              �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?�������?�q�q�?9��8���?              �?�������?333333�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?      �?              �?      �?        �m۶m��?%I�$I��?      �?      �?F]t�E�?]t�E]�?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        (�����?�k(���?      �?                      �?��hgJ��?��%f-�?�.�袋�?F]t�E�?      �?        �������?�������?�������?�������?      �?                      �?      �?        Y]����?�rS�<�v?      �?        ��7��M�?d!Y�B�?�?�?      �?      �?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���bhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKՅ�h��B@5         .                   �c@��Wޫ��?�           ��@               )                    �?p=
ף0�?_             d@                     	          �����fv�S��?6            �T@        ������������������������       �                     @                                   �?���B���?4            �S@                                   �C@�q�����?             9@        ������������������������       �                      @               	                    �?\X��t�?             7@        ������������������������       �                     �?        
              
             �?�eP*L��?             6@                     
             �?���|���?	             &@        ������������������������       �                     �?                                  �c@�z�G��?             $@                                 @_@      �?              @                                  �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                   �?���!pc�?             &@        ������������������������       �                     �?                                  �d@z�G�z�?             $@                                 @_@�����H�?             "@                                  �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               (                    @N@�&=�w��?             �J@              #       
             �?�>����?             ;@                      	          033�?���7�?             6@        ������������������������       �                     (@        !       "                   �`@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        $       '                   a@z�G�z�?             @        %       &                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        *       +       	          033@ ���J��?)            �S@       ������������������������       �        '            �R@        ,       -       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        /       �                    �?�i禺h�?u           ��@       0       i       
             �?��,���?�            �v@        1       B                   P`@���N��?M             ]@        2       7                     L@�'�`d�?            �@@        3       6                     F@�C��2(�?	             &@        4       5                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        8       9       	          ����?���!pc�?             6@        ������������������������       �                     @        :       =                    @M@ҳ�wY;�?             1@        ;       <       	             �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        >       ?                    `P@�C��2(�?             &@       ������������������������       �                      @        @       A                   �[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        C       `                   @q@F~��7�?6            �T@       D       O                    @L@҄��?+            �P@       E       F                    �?z�G�z�?             D@        ������������������������       �                     2@        G       N       	             @�X����?             6@       H       I                    �?      �?             4@        ������������������������       �                     @        J       K                   �`@�t����?             1@       ������������������������       �        	             ,@        L       M       	          @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        P       Y                   �l@�n_Y�K�?             :@       Q       R                   p`@�E��ӭ�?             2@        ������������������������       �                      @        S       X                   �d@     ��?
             0@       T       W                   h@@4և���?	             ,@        U       V                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        Z       [       
             �?      �?              @        ������������������������       �                     �?        \       _                   �n@և���X�?             @       ]       ^       	          ���@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        a       h                    �?�t����?             1@       b       g                   �c@X�Cc�?             ,@        c       d                     J@����X�?             @        ������������������������       �                     @        e       f                    �M@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        j       w                    @L@��GEI_�?�            �n@       k       p                    �?@�E�x�?|            �h@        l       o                    @F@r�q��?             2@        m       n       	          ����?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             (@        q       v                    \@@~��?o            @f@        r       s                    �I@      �?             @@       ������������������������       �                     8@        t       u                   �[@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        Y            @b@        x       {                    �?      �?             H@        y       z                   �b@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        |       �       	          033@�MI8d�?            �B@       }       �                    �?l��\��?             A@        ~       �                     N@      �?              @               �                    �?      �?             @       �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        ������������������������       �                     @        �       �                    �?�8l�9��?�            �j@       �       �       	          033�?*
;&���?}             g@        �       �                   �s@j���� �?             A@       �       �                    _@8^s]e�?             =@        ������������������������       �                     @        �       �       	          833�?�û��|�?             7@       �       �                    �?�E��ӭ�?             2@        ������������������������       �                     @        �       �                    �N@�q�q�?
             (@       �       �                   `Z@      �?              @        ������������������������       �                     �?        �       �                   Pg@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       �       �                    @K@z�G�z�?             @        �       �                   `m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          hff�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Lͩ�?c            �b@       �       �                     E@�X�C�?M             \@        �       �                    b@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?0��_��?I            �Z@       �       �       
             �?XI�~�?9            @S@        ������������������������       �                     $@        �       �                   �j@t�e�í�?2            �P@        �       �       	             �?r�q��?             2@        �       �                   i@�q�q�?             @        ������������������������       �                      @        �       �                   @_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @b@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �s@@9G��?'            �H@       �       �                    c@ qP��B�?#            �E@       ������������������������       �                      D@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �t@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `\@д>��C�?             =@        �       �       	             @����X�?             @       �       �                   �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        �       �       	          033�?P�Lt�<�?             C@       ������������������������       �                     6@        �       �                   @^@      �?
             0@        �       �                   �c@z�G�z�?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �       	          ���@      �?             >@       �       �                   �`@���Q��?             9@       �       �                   �[@���y4F�?             3@        �       �                    �O@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  +^�ɑA�?�P47��?�������?�������?�]�ڕ��?��]�ڕ�?      �?        ى�؉��?��؉���?�p=
ף�?���Q��?              �?!Y�B�?��Moz��?      �?        t�E]t�?]t�E�?F]t�E�?]t�E]�?      �?        333333�?ffffff�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        F]t�E�?t�E]t�?              �?�������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�x+�R�?tHM0���?h/�����?�Kh/��?F]t�E�?�.�袋�?              �?�������?�������?              �?      �?        �������?�������?      �?      �?      �?                      �?              �?              �?�A�A�?��-��-�?              �?      �?      �?      �?                      �?)�k�,�?�#(ͦ�?}�'}�'�?�`�`�?j��FX�?�=�����?'�l��&�?6�d�M6�?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?t�E]t�?F]t�E�?              �?�������?�������?�������?UUUUUU�?      �?                      �?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?      �?        ���ˊ��?��h���?�d�M6��?N6�d�M�?ffffff�?ffffff�?      �?        �E]t��?]t�E]�?      �?      �?              �?<<<<<<�?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?ى�؉��?;�;��?r�q��?�q�q�?      �?              �?      �?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?�������?�������?�m۶m��?%I�$I��?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?                      �?              �?�d����?;ڼOqɰ?և���X�?9/���?�������?UUUUUU�?      �?      �?              �?      �?              �?        ��G?���?p�\�w?      �?      �?      �?              �?      �?      �?                      �?      �?              �?      �?]t�E�?t�E]t�?      �?                      �?��L���?L�Ϻ��?------�?�������?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?              �?                      �?�ީk9��?`����?8��Moz�?���,d!�?ZZZZZZ�?�������?	�=����?|a���?              �?��,d!�?8��Moz�?r�q��?�q�q�?              �?�������?�������?      �?      �?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?�������?�������?      �?      �?      �?                      �?      �?              �?                      �?�������?�������?      �?                      �?      �?        �K~��?�6�i�?n۶m۶�?�$I�$I�?      �?      �?              �?      �?        �V�9�&�?"5�x+��?V~B����?5�wL��?              �?�rv��?�1����?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        9/���?������?�}A_З?��}A�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?UUUUUU�?�������?      �?                      �?|a���?a���{�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?(�����?���k(�?              �?      �?      �?�������?�������?              �?      �?      �?      �?                      �?              �?      �?      �?333333�?�������?6��P^C�?(������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ+�MhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKх�h��B@4         �       
             �?.��X~��?�           ��@                                 �a@�+$�jP�?            {@                      
             �?0�)AU��?E            �\@                      	          033�?��S�ۿ?	             .@                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        	       
                   �c@`�LVXz�?<            �X@       ������������������������       �        0            @S@                                   �P@���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?               A                    �?�c�����?�            �s@               8       	          033�?N1���?Q            �^@                                  �?X�<ݚ�?:            �V@                      	          ����?<���D�?            �@@                                  �?������?             .@                                 `j@      �?              @        ������������������������       �                      @                                  �[@�q�q�?             @        ������������������������       �                     �?                                   �?z�G�z�?             @        ������������������������       �                     @                                   @J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@               #       	          ����?p�ݯ��?&            �L@                                   �d@���7�?             6@       ������������������������       �        
             3@        !       "       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        $       )                   �^@և���X�?            �A@        %       (                    �?$�q-�?             *@        &       '                   `]@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        *       7                   xr@���|���?             6@       +       4                   �`@�d�����?             3@        ,       /                    �?      �?              @        -       .                   �m@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        0       3                    `@      �?             @        1       2                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        5       6       	          833�?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        9       @                   �e@     ��?             @@       :       ?                   d@�r����?             >@       ;       <                    @@4և���?             <@       ������������������������       �                     9@        =       >                   0`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        B       O                    �?�+�$f��?~            �h@        C       L                   �b@      �?             <@       D       E                   `a@�LQ�1	�?             7@        ������������������������       �                     &@        F       K                    �L@      �?             (@        G       H                   �b@���Q��?             @        ������������������������       �                      @        I       J                   u@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        M       N                     L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        P       s       	          ����?4և����?k             e@        Q       h                    �?�x
�2�?2            �R@       R       [                    @G@ܷ��?��?(             M@        S       V                   �\@�q�q�?             "@        T       U                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        W       X       	          ����?r�q��?             @        ������������������������       �                     @        Y       Z                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        \       a       	          `ff�?��<D�m�?!            �H@        ]       `                    \@z�G�z�?             $@        ^       _       	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        b       c                   `_@ ���J��?            �C@       ������������������������       �                     :@        d       g                   Pi@$�q-�?	             *@        e       f                   i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        i       p                    �?     ��?
             0@       j       m       	          033�?�	j*D�?             *@       k       l                   @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        n       o                   �b@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        q       r                    ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        t       {                   �j@`�q�0ܴ?9            �W@        u       v       	          `ff�?�����H�?             2@        ������������������������       �                     �?        w       z                    �H@�IєX�?             1@        x       y                   h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        |       }                    @M@P�Lt�<�?-             S@       ������������������������       �                    �B@        ~                           c@�7��?            �C@       ������������������������       �                    �B@        ������������������������       �                      @        �       �                    �K@h������?�            �r@       �       �                   Pd@���Lͩ�?�             l@       �       �       	            �?,�� ��?�            �k@       �       �                    �?Hx�i�.�?o             g@        �       �                    `@:	��ʵ�?            �F@       �       �                   pb@�ՙ/�?             5@        ������������������������       �                     "@        �       �                   �c@�q�q�?             (@        ������������������������       �                     @        �       �                   Pl@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �        V            �a@        �       �                    �?<ݚ)�?             B@        ������������������������       �                     0@        �       �       	             �?�G�z��?             4@       �       �                    �?����X�?             ,@       �       �                    �J@z�G�z�?             $@       �       �       	             �?      �?              @        ������������������������       �                     @        �       �                    �F@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   e@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?rOP\6�?7            @S@       �       �                    �?�G�z��?             D@       �       �                    �?�P�*�?             ?@        �       �                    �M@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?�q�q�?             5@       �       �                    �?��
ц��?
             *@        ������������������������       �                     @        �       �                   `l@���Q��?             $@       �       �                    @O@      �?              @       �       �                    �?z�G�z�?             @       �       �                     M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �m@      �?              @       ������������������������       �                     @        �       �                    @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?��G���?            �B@        �       �                    �M@��S�ۿ?
             .@        �       �                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                    �P@���!pc�?             6@       �       �       	             @      �?             0@       �       �                   �a@�θ�?
             *@        ������������������������       �                     @        �       �                   �_@      �?             @        ������������������������       �                     �?        �       �       	          ����?���Q��?             @       �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  ��� ���?���o���?B{	�%��?/�����?p�}��?��Gp�?�?�������?      �?      �?              �?      �?                      �?[�R�֯�?�~�@��?              �?F]t�E�?�.�袋�?              �?      �?        :�&oe�?�V�9�&�?�}�K�`�?�:ڼO�?r�q��?�q�q�?|���?|���?wwwwww�?�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?      �?                      �?      �?              �?        Cy�5��?^Cy�5�?F]t�E�?�.�袋�?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?�؉�؉�?;�;��?�������?UUUUUU�?              �?      �?              �?        F]t�E�?]t�E]�?y�5���?Cy�5��?      �?      �?      �?      �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?        F]t�E�?]t�E�?      �?                      �?      �?              �?      �?�?�������?�$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        /�����?�Cc}h�?      �?      �?Y�B��?��Moz��?              �?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?                      �?�m۶m۶?I�$I�$�?o0E>��?�n0E>�?a���{�?��=���?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?և���X�?��S�r
�?�������?�������?      �?      �?              �?      �?                      �?�A�A�?��-��-�?              �?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?      �?;�;��?vb'vb'�?      �?      �?      �?                      �?333333�?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?W�+�ɥ?��F}g��?�q�q�?�q�q�?      �?        �?�?      �?      �?              �?      �?                      �?(�����?���k(�?              �?�A�A�?��[��[�?              �?      �?        ��jg���?��Tb*1�?�6�i�?�K~��?ݵ?ݵ?�?QQ�?��X���?@bw�#�?��O��O�?l�l��?�<��<��?�a�a�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��8��8�?�8��8��?      �?        �������?�������?�$I�$I�?�m۶m��?�������?�������?      �?      �?              �?      �?      �?      �?                      �?      �?      �?              �?      �?              �?      �?              �?      �?        �������?UUUUUU�?      �?                      �?      �?      �?              �?      �?        ��O����?dj`��?�������?�������?�RJ)���?�Zk����?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?�;�;�?�؉�؉�?      �?        �������?333333�?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?      �?      �?      �?              �?      �?      �?                      �?              �?#�u�)��?v�)�Y7�?�������?�?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?t�E]t�?      �?      �?ى�؉��?�؉�؉�?      �?              �?      �?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJY]hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKǅ�h��B�1         �       
             �?��;/M�?�           ��@                                 0b@@�0�!��?           �{@                                   �?���1��?B            �Z@       ������������������������       �        4            �T@               
                    �? �q�q�?             8@               	                    �?؇���X�?             @                                   @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             1@               /                    �?�Ks1���?�            �t@               .                   `c@      �?/             S@              '                    �?�G\�c�?(            @P@                                  �?b�2�tk�?             B@                      	          ����?���Q��?	             .@        ������������������������       �                     @                                   �M@      �?              @                                   `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �N@r�q��?             @        ������������������������       �                     @                                  Xs@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �e@���N8�?             5@        ������������������������       �                     �?               &       	          ����?z�G�z�?             4@               #                   �p@      �?              @               "                    @N@      �?             @               !                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        $       %                   �t@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             (@        (       )                   `X@д>��C�?             =@        ������������������������       �                      @        *       -                    �?�����H�?             ;@        +       ,                   @q@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             0@        ������������������������       �                     &@        0       y       	          ����?��L~1_�?�            0p@       1       `                   �n@�rF���?j            �d@       2       I                    �?�j&|mH�?=            @X@        3       :       	          ����?�e����?            �C@        4       5       
             �?���y4F�?             3@        ������������������������       �                     �?        6       9                    �E@r�q��?             2@        7       8                    �C@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ;       H                   �c@���Q��?             4@       <       =                    �G@��.k���?             1@        ������������������������       �                     @        >       ?                    `@և���X�?
             ,@        ������������������������       �                     @        @       A       	          ����?�eP*L��?             &@        ������������������������       �                     @        B       C                   `_@r�q��?             @        ������������������������       �                     @        D       E                   �k@�q�q�?             @        ������������������������       �                     �?        F       G                    m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        J       Q                   `_@V�a�� �?$             M@        K       P                   j@@4և���?             <@        L       M                    �K@����X�?             @        ������������������������       �                     @        N       O                    �M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        R       _                   �m@�q�q�?             >@       S       ^                    �?����X�?             <@       T       U       	          ����?X�<ݚ�?             2@        ������������������������       �                     @        V       W                   �\@�n_Y�K�?             *@        ������������������������       �                     @        X       ]                    �?����X�?             @       Y       Z                   �_@�q�q�?             @        ������������������������       �                      @        [       \                   �`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        a       p                    �?�t����?-             Q@       b       o                   �e@�:�]��?!            �I@       c       h                    �? "��u�?              I@        d       g                   @^@�t����?             1@        e       f                   (r@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        i       n                    `@Pa�	�?            �@@        j       m       	          433�?z�G�z�?             @        k       l                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        ������������������������       �                     �?        q       x                    �?������?             1@       r       w                   �s@�q�q�?	             (@       s       v                   �_@�����H�?             "@        t       u       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        z       {                   �Z@��V�I��?<            �W@        ������������������������       �                     �?        |       }                   �p@����D��?;            @W@       ������������������������       �        +            @Q@        ~       �                    `Q@�8��8��?             8@              �                   �e@�nkK�?             7@       ������������������������       �                     5@        �       �       	          ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�&����?�            @r@       �       �                     L@��2(&�?�            @n@       �       �       	             @PÅ�R1�?}            �f@       �       �                    c@�ȨF=�?|            `f@        �       �                   �`@      �?              @        �       �                   �R@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �A@`RI��d�?w            `e@        �       �                   �c@@4և���?             ,@        �       �                   pc@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�#��g1�?k            �c@        �       �                    �?l��\��?             A@       �       �       	            �?`Jj��?             ?@       �       �                    �I@ 7���B�?             ;@       ������������������������       �                     5@        �       �                   @_@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          hff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        R            �^@        ������������������������       �                      @        �       �                    �?�u���?&            �N@        �       �                    s@ףp=
�?             4@       ������������������������       �                     (@        �       �                    �?      �?              @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?D^��#��?            �D@        �       �                    �P@�q�q�?             5@       �       �                   d@������?
             1@       ������������������������       �                     *@        ������������������������       �                     @        �       �                   0b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �M@      �?             4@        ������������������������       �                     &@        �       �                   �]@X�<ݚ�?	             "@        ������������������������       �                      @        �       �                    �?����X�?             @        �       �                   �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@`�Q��?              I@        �       �                    \@������?             1@        ������������������������       �                     "@        �       �                    @K@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �U@�C��2(�?            �@@        ������������������������       �                     @        ������������������������       �                     >@        �t�b�@     h�h)h,K ��h.��R�(KK�KK��hb�Bp  �X�5��?�S�$e�?�������?ZZZZZZ�?�+J�#�?�S�rp��?              �?UUUUUU�?�������?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?              �?��Ͽk�?�:��?      �?      �?S+�R+��?[��Z���?9��8���?�8��8��?333333�?�������?      �?              �?      �?      �?      �?      �?                      �?UUUUUU�?�������?              �?      �?      �?              �?      �?        ��y��y�?�a�a�?      �?        �������?�������?      �?      �?      �?      �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?              �?a���{�?|a���?              �?�q�q�?�q�q�?F]t�E�?t�E]t�?      �?                      �?      �?                      �?c4�w-F�?��t.�?�־a��?yJ���?���fy�?w�<�L��?�A�A�?�-��-��?(������?6��P^C�?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?333333�?�������?�������?�?      �?        ۶m۶m�?�$I�$I�?              �?t�E]t�?]t�E�?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        a���{�?��{a�?�$I�$I�?n۶m۶�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?�q�q�?r�q��?              �?;�;��?ى�؉��?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?              �?      �?        �?<<<<<<�?�?}}}}}}�?���Q��?�G�z�?�?<<<<<<�?�$I�$I�?�m۶m��?              �?      �?                      �?|���?|���?�������?�������?      �?      �?      �?                      �?              �?              �?      �?        �?xxxxxx�?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?      �?      �?                      �?              �?      �?                      �?AL� &W�?<�����?      �?        X`��?P?���O�?              �?UUUUUU�?UUUUUU�?d!Y�B�?�Mozӛ�?              �?      �?      �?              �?      �?              �?        *T�P��?�W�^�z�?��.���?t�E]t�?�!H��h�?��}kdu�?�R"x���?���}��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?��_@�?@���?n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?        >"'wc�?A����?------�?�������?���{��?�B!��?	�%����?h/�����?      �?        �������?UUUUUU�?              �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?T\2�h�?XG��).�?�������?�������?      �?              �?      �?      �?      �?              �?      �?              �?        �]�ڕ��?,Q��+�?UUUUUU�?UUUUUU�?xxxxxx�?�?      �?                      �?      �?      �?              �?      �?              �?      �?              �?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        ��(\���?{�G�z�?�?xxxxxx�?              �?      �?      �?      �?                      �?]t�E�?F]t�E�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ4
hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK݅�h��B@7         ~       
             �?���:���?�           ��@              +                   a@lRV����?�            �x@                                  �?���m��?�            �n@                      	          pff�?��>4և�?             <@                      	          @33�?      �?	             0@        ������������������������       �                     �?                                   d@��S�ۿ?             .@       ������������������������       �                     &@        	       
                    �L@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                    P@      �?	             (@       ������������������������       �                     "@        ������������������������       �                     @               "       	          ����?���s�?�             k@               !                   �[@��`qM|�?4            �T@                                  �L@�ʈD��?            �E@                                   �?�S����?             3@                     	             �?�����H�?             2@       ������������������������       �                     (@                                  o@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                    �? �q�q�?             8@                                  �?@4և���?             ,@                     	          ����?ףp=
�?             $@        ������������������������       �                     @                                  �Y@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     D@        #       *                    �D@ 
�V�?Y            �`@        $       )                    �?z�G�z�?             @       %       &                     C@      �?             @        ������������������������       �                      @        '       (                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        U             `@        ,       ;                    �G@���}��?`             c@        -       0                    �?��%��?            �B@        .       /                    Z@@4և���?	             ,@        ������������������������       �                     �?        ������������������������       �                     *@        1       8                    �?8����?             7@       2       3                   �Z@r�q��?	             2@        ������������������������       �                     �?        4       5                    �E@�t����?             1@       ������������������������       �                     ,@        6       7                    b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        9       :                     D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        <       I                   �_@z�G�z�?K            �\@        =       >                   �h@����X�?             <@        ������������������������       �                     "@        ?       @                    �H@D�n�3�?             3@        ������������������������       �                     @        A       D                   @]@��S���?             .@        B       C       	          `ff�?      �?              @        ������������������������       �                      @        ������������������������       �                     @        E       F       	             �?؇���X�?             @       ������������������������       �                     @        G       H                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        J       K                   0a@д>��C�?8            �U@        ������������������������       �                     �?        L       _                    �?�T|n�q�?7            �U@        M       T                    �J@����X�?             5@        N       O                    �?      �?              @        ������������������������       �                      @        P       Q                   �`@�q�q�?             @        ������������������������       �                     @        R       S                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        U       ^                    �?8�Z$���?             *@       V       ]                    �?      �?              @       W       \                    @O@؇���X�?             @       X       [                   �c@      �?             @        Y       Z                   Xs@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        `       m                    �?�?�<��?(            @P@       a       b                     L@������?            �D@        ������������������������       �                     3@        c       d                   @a@�C��2(�?             6@        ������������������������       �                     &@        e       f                   �f@"pc�
�?             &@        ������������������������       �                     @        g       h                   h@����X�?             @        ������������������������       �                     �?        i       l                   �a@r�q��?             @        j       k       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        n       {                    �?      �?             8@       o       v                    �N@z�G�z�?             4@       p       q       	          ����?      �?	             0@        ������������������������       �                     &@        r       u                   �`@z�G�z�?             @        s       t                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        w       z                    @      �?             @       x       y                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        |       }                   �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @               �                    _@Mm7�?�            u@        �       �                    @K@8�A�0��?              F@        �       �                    �?R���Q�?             4@       �       �                   `V@�X�<ݺ?             2@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                      @        �       �       	          ����?      �?             8@       �       �                   �`@�	j*D�?
             *@       ������������������������       �                     @        �       �                    �N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        �       �                    �?��S�U�?�            Pr@       �       �                   @E@���ZG�?�            p@        �       �                   �a@���Q��?             $@        ������������������������       �                     @        �       �       	          @33�?؇���X�?             @        �       �                    �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             @أ����?�            �n@       �       �                   �`@� �$m�?�            �n@       �       �                    �?4/Gjϵ?a            �c@       �       �                   pc@P���Q�?W            �a@        �       �       	            �?     ��?(             P@       ������������������������       �        "            �J@        �       �                    �?�C��2(�?             &@        ������������������������       �                      @        �       �                   @n@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����?�˹�m��?/             S@       �       �                    �?Hn�.P��?%             O@        �       �                   `\@�θ�?             *@        ������������������������       �                      @        �       �                    �?�C��2(�?             &@       �       �                   �d@؇���X�?             @        ������������������������       �                     @        �       �                   pr@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �H@        �       �                    �?d}h���?
             ,@        �       �       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             1@        �       �                    �?      �?2             V@       �       �                    �K@$��$�L�?-            �S@       ������������������������       �                     I@        �       �       	          @33�?�c�Α�?             =@       �       �                   �m@��S���?	             .@        ������������������������       �                     @        �       �                    �?���!pc�?             &@        �       �                    �N@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    k@@4և���?             ,@        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        �       �       	          833�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �r@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    f@      �?             B@       �       �                    k@�P�*�?             ?@        �       �                    �?�8��8��?	             (@       ������������������������       �                     @        �       �                   `b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?p�ݯ��?             3@       �       �                    a@���|���?             &@        ������������������������       �                      @        �       �                     L@�<ݚ�?             "@       ������������������������       �                     @        �       �       	          @33�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  !��Q��?p��1W-�?O�+�	��?�	�����?򸳄���?�iOd �?۶m۶m�?I�$I�$�?      �?      �?              �?�������?�?      �?              �?      �?      �?                      �?      �?      �?              �?      �?        �`^0/��?�}�>C�?��k���?�@	o4u�?�}A_з?A_���?^Cy�5�?(������?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?�$I�$I�?n۶m۶�?�������?�������?              �?�������?�������?              �?      �?                      �?              �?              �?g��1�~?������?�������?�������?      �?      �?              �?      �?      �?              �?      �?                      �?              �?������?(������?���L�?}���g�?n۶m۶�?�$I�$I�?              �?      �?        8��Moz�?d!Y�B�?UUUUUU�?�������?      �?        �?<<<<<<�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?�������?�������?�$I�$I�?�m۶m��?              �?(������?l(�����?              �?�?�������?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?|a���?a���{�?      �?        6eMYS��?���)k��?�$I�$I�?�m۶m��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?      �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?              �?      �?                      �? �����?�����?������?p>�cp�?              �?F]t�E�?]t�E�?              �?F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?      �?�������?�������?      �?      �?              �?�������?�������?      �?      �?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?������?�Ed����?颋.���?/�袋.�?333333�?333333�?��8��8�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?vb'vb'�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�� S�1�?P����8�?=�<�<��?���?�������?333333�?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?���h�?�KA���?еʆ#��?�Q���β?�O[h���?�Kz�Ӧ?ffffff�?�������?     ��?      �?      �?        ]t�E�?F]t�E�?      �?        �q�q�?�q�q�?      �?                      �?��P^Cy�?^Cy�5�?t�9�s�?�c�1ƨ?ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?              �?        I�$I�$�?۶m۶m�?      �?      �?              �?      �?              �?              �?              �?      �?��]-n��?�3���?      �?        5�rO#,�?�{a���?�?�������?              �?F]t�E�?t�E]t�?333333�?�������?              �?      �?        �������?UUUUUU�?      �?                      �?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?�Zk����?�RJ)���?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?              �?      �?        ^Cy�5�?Cy�5��?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?              �?      �?      �?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��;hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKم�h��B@6         �       	          ����?({E�B��?�           ��@              W       
             �?�*�?(           �}@                                  �e@vp�*�?�             h@                                  �O@ �й���?0            @R@                                  �?@	tbA@�?,            @Q@                      	          ����?��?^�k�?            �A@                                 `X@ ��WV�?             :@               	                    �?      �?              @       ������������������������       �                     @        
                           �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     "@        ������������������������       �                     A@        ������������������������       �                     @               @                   `a@��Q��?R             ^@                                 �]@
j*D>�?4            �S@                      	          ����?؇���X�?             5@       ������������������������       �                     ,@                                    L@և���X�?             @                                  �?z�G�z�?             @        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @               ?                   �`@�\��N��?&            �L@              0                   `b@     ��?!             H@              /                    �?X�Cc�?             <@                                   @C@��<b���?             7@        ������������������������       �                     �?        !       .                   �`@"pc�
�?             6@       "       )                    �M@؇���X�?             5@       #       (                   �a@�IєX�?             1@       $       %                    �?�����H�?             "@       ������������������������       �                     @        &       '                   0l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        *       +                    @N@      �?             @        ������������������������       �                     �?        ,       -       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        1       >                    �N@R���Q�?             4@       2       =                    �?�KM�]�?             3@       3       6                   �k@r�q��?
             (@        4       5                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        7       8                   @d@ףp=
�?             $@        ������������������������       �                     @        9       :                    @J@      �?             @        ������������������������       �                      @        ;       <                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        A       F                   `_@d}h���?             E@        B       E                    m@�X�<ݺ?             2@        C       D                    b@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        G       L                   p`@�q�q�?             8@        H       I                    �?����X�?             @        ������������������������       �                     @        J       K                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        M       N                     L@@�0�!��?             1@        ������������������������       �                     @        O       P                   0h@�z�G��?             $@        ������������������������       �                      @        Q       R                    �?      �?              @        ������������������������       �                     @        S       T                    �?      �?             @        ������������������������       �                      @        U       V                     P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        X                           �? ��z��?�            �q@       Y       `                   �e@     ��?�             p@        Z       [                    �?����X�?             <@        ������������������������       �                     @        \       ]       	          833�?r�q��?             8@       ������������������������       �                     1@        ^       _                   ``@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        a       n                     L@p�|�i�?�            �l@       b       m                    �?�Y�ߠ?i            `f@        c       h                    @F@t��ճC�?             F@        d       e                   �p@؇���X�?             ,@        ������������������������       �                      @        f       g                   pc@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        i       j                   �c@(;L]n�?             >@       ������������������������       �                     8@        k       l                   `\@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        Q            �`@        o       ~                     P@�q��/��?            �H@       p       {                    b@b�h�d.�?            �A@       q       z                    �?      �?             @@       r       u                   0b@r�q��?             8@        s       t       	          @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        v       w                   `a@�����?             5@       ������������������������       �                     &@        x       y                    �O@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        |       }                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   �Y@|��?���?             ;@        ������������������������       �                     $@        �       �                    �?������?             1@       �       �                    @P@      �?              @       �       �                   `_@�q�q�?             @        ������������������������       �                     �?        �       �                   Pn@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?�T|n�q�?�             p@        �       �                   �b@���=A�?4             S@       �       �       	          ��� @^l��[B�?)             M@       �       �                    �?P����?             C@        �       �                   `Y@�n_Y�K�?             *@        ������������������������       �                     @        �       �       
             �?z�G�z�?             $@       �       �                   �Z@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       	             �?z�G�z�?             9@        ������������������������       �                     @        �       �                    �?�C��2(�?             6@       �       �                   �k@�X�<ݺ?             2@       ������������������������       �        	             (@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        �       �                    �?�q�q�?             2@       �       �                    �?      �?              @        ������������������������       �                     @        �       �                   Pd@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        �       �       	          ����?�h�ഭ�?i            �f@        �       �                    �G@�חF�P�?"             O@        �       �       
             �?z�G�z�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�KM�]�?            �L@       �       �                   @_@��<D�m�?            �H@       ������������������������       �                    �@@        �       �                    ^@     ��?	             0@        ������������������������       �                      @        �       �                   P`@@4և���?             ,@       ������������������������       �                     &@        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        �       �                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �O@      �?              @       �       �                   �`@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�S���?G             ^@       �       �                    �?,���$�?6            @X@       �       �                   `b@������?2            @V@       �       �       
             �?P�Lt�<�?,             S@       �       �                     R@�k~X��?(             R@       ������������������������       �        '            �Q@        ������������������������       �                     �?        �       �                   `W@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �]@�n_Y�K�?             *@        ������������������������       �                      @        �       �                    �?���!pc�?             &@        ������������������������       �                     @        �       �       	          ����?և���X�?             @        ������������������������       �                     @        �       �                    �L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     7@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  Ac�Zb�?`yΨ�N�?��ԋ���?�V�V�?c�z���?�~����?����?����Ǐ�?ہ�v`��?�%~F��?�A�A�?_�_��?;�;��?O��N���?      �?      �?              �?      �?      �?      �?                      �?              �?              �?              �?              �?ffffff�?�������?;�;��?b'vb'v�?�$I�$I�?۶m۶m�?              �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?      �?      �?                      �?      �?        y�5���?�5��P�?      �?      �?%I�$I��?�m۶m��?��,d!�?��Moz��?              �?/�袋.�?F]t�E�?۶m۶m�?�$I�$I�?�?�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?333333�?333333�?(�����?�k(���?UUUUUU�?�������?      �?      �?              �?      �?        �������?�������?              �?      �?      �?              �?      �?      �?              �?      �?                      �?      �?              �?        ۶m۶m�?I�$I�$�?�q�q�?��8��8�?UUUUUU�?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?�������?ZZZZZZ�?              �?333333�?ffffff�?      �?              �?      �?              �?      �?      �?              �?      �?      �?      �?                      �?ǬӢ�~�?șb��
�?     ��?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        �k(����?^Cy�5�?�l|3�v�?�ir�y)�?�E]t��?t�E]t�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�?      �?        �������?UUUUUU�?              �?      �?              �?        /����?և���X�?;��:���?_�_��?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?=��<���?�a�a�?      �?        �������?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        	�%����?{	�%���?              �?xxxxxx�?�?      �?      �?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        6eMYS��?���)k��?�P^Cy�?��P^Cy�?��=���?�=�����?Q^Cy��?�P^Cy�?;�;��?ى�؉��?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?      �?        F]t�E�?]t�E�?�q�q�?��8��8�?              �?UUUUUU�?�������?              �?      �?              �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?              �?      �?              �?        �~�~�?-�-��?��RJ)��?�Zk����?�������?�������?      �?      �?      �?                      �?      �?        (�����?�k(���?և���X�?��S�r
�?              �?      �?      �?      �?        �$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?�$I�$I�?�m۶m��?              �?      �?              �?        �����ݭ?""""""�?���fy�?�,O"Ӱ�?B�P�"�?ؽ�u�{�?(�����?���k(�?�q�q�?�8��8��?              �?      �?              �?      �?      �?      �?      �?                      �?              �?ى�؉��?;�;��?      �?        t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?              �?      �?      �?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJS�)/hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK˅�h��B�2         �       
             �?��}���?�           ��@              =                    �?�����?           �y@                                   �?����r��?h            �c@                                  @L@�$�����?8            @T@                                  `p@���N8�?             E@       ������������������������       �                    �@@                                  �`@�<ݚ�?             "@              	                    �D@���Q��?             @        ������������������������       �                      @        
                           �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                  �r@x�����?            �C@                                  �?l��\��?             A@                                   �?@�0�!��?             1@                                  �?��S�ۿ?
             .@                                  �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     @               6                    �?v�(��O�?0            �R@                                  ]@L
�q��?&            �M@                                  @e@�z�G��?             $@       ������������������������       �                     @                      	          @33�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                3                   @b@�D��?            �H@       !       2                   �`@��r._�?            �D@       "       /                    @>���Rp�?             =@       #       &       	          ����?z�G�z�?             9@        $       %                    @L@      �?             @        ������������������������       �                      @        ������������������������       �                      @        '       ,       	          `ff�?؇���X�?             5@       (       )                   �b@�IєX�?
             1@       ������������������������       �                     &@        *       +                    �K@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        -       .                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        0       1                   �r@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        4       5       	          ����?      �?              @       ������������������������       �                     @        ������������������������       �                      @        7       <                   8r@      �?
             0@       8       9                   `b@z�G�z�?	             .@       ������������������������       �                     &@        :       ;                   �`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        >       }                   �b@0����?�            �o@       ?       H                   i@|�U�7��?�             n@        @       A                    �?`׀�:M�?-            �R@       ������������������������       �        !             L@        B       G                    �N@�X�<ݺ?             2@        C       D                    �M@�����H�?             "@       ������������������������       �                     @        E       F                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        I       L                   �Z@�A�D6h�?p            �d@        J       K       	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        M       Z                    �?|E+�	��?m            @d@        N       O                    �?ȵHPS!�?             :@        ������������������������       �                     @        P       Q       	             �?�S����?             3@        ������������������������       �                     @        R       Y                   �b@z�G�z�?	             .@       S       T                   �j@���!pc�?             &@        ������������������������       �                     @        U       V                    �?      �?             @        ������������������������       �                      @        W       X                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        [       |                   0a@����p�?^             a@       \       o       	          ����?�H�@=��?M            �[@        ]       ^                   Pi@PN��T'�?&             K@        ������������������������       �                     @        _       n       	          ����?`�H�/��?%            �I@       `       m                   �`@�חF�P�?             ?@       a       b                    @K@�r����?             >@        ������������������������       �        	             1@        c       h                    \@�	j*D�?             *@        d       e                   @_@      �?             @        ������������������������       �                      @        f       g                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        i       l                   �`@؇���X�?             @        j       k                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        p       y                    �R@���U�?'            �L@       q       x                   xp@ �Jj�G�?%            �K@       r       s       
             �?h�����?             <@        ������������������������       �                     @        t       u                   8p@�nkK�?             7@       ������������������������       �                     5@        v       w                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ;@        z       {                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@        ~       �                   Pc@      �?	             (@              �                    �D@      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @       �       �                     K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��=��?�            Pt@        �       �       	          ����?�0���8�?C            @[@       �       �                   �b@�G�5��?(            @Q@       �       �                   �j@�X�<ݺ?             B@        �       �                    �?�t����?
             1@       �       �                    �?      �?	             0@        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     3@        �       �                    �I@�eP*L��?            �@@        �       �       	          ����?�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        �       �                   `a@���Q��?             4@       �       �                   pk@��
ц��?             *@        ������������������������       �                     @        �       �                   �e@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                    @O@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @b@��Q���?             D@       �       �                    �?؇���X�?             <@        �       �       	          `ff�?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                    @N@���}<S�?             7@       �       �                   �`@�r����?             .@        ������������������������       �                     @        �       �                   �`@      �?              @        ������������������������       �                     �?        �       �                    �J@؇���X�?             @        ������������������������       �                     @        �       �                    @K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             (@       �       �                    �?      �?              @       ������������������������       �                     @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ���@p)�����?�             k@       �       �                   �c@(;L]n�?�            @j@       �       �                   �^@io8�?H             ]@        �       �                    �?����?�?            �F@        �       �                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     E@        �       �                    _@@�j;��?-            �Q@        ������������������������       �                     @        �       �                   �c@ =[y��?,             Q@       �       �                   �s@ ����?*            @P@       ������������������������       �        '             N@        �       �                   (t@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        :            �W@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  q��H��?��>���?�Q�c	�?������?�[��[��?� � �?X�<ݚ�?uk~X��?�a�a�?��y��y�?              �?�q�q�?9��8���?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�A�A�?��o��o�?�������?------�?�������?ZZZZZZ�?�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?      �?        Y�%�X�?O贁N�?��V'�?�pR���?333333�?ffffff�?              �?      �?      �?              �?      �?        ������??4և���?�ڕ�]��?ە�]���?�i��F�?GX�i���?�������?�������?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?�?�?      �?        �������?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?      �?              �?      �?              �?              �?      �?              �?      �?              �?      �?�������?�������?              �?      �?      �?      �?                      �?      �?        '���H�?[
����?���?>&�=&��?к����?��L��?              �?�q�q�?��8��8�?�q�q�?�q�q�?              �?      �?      �?              �?      �?                      �?Nk�OT�?�2	v��?�������?�������?              �?      �?        �n���??,R�n�?�؉�؉�?��N��N�?              �?^Cy�5�?(������?              �?�������?�������?t�E]t�?F]t�E�?              �?      �?      �?      �?              �?      �?      �?                      �?              �?�����Ҳ?�������?q��$�?��+c��?h/�����?&���^B�?      �?        �?�������?��RJ)��?�Zk����?�?�������?              �?;�;��?vb'vb'�?      �?      �?              �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?                      �?p�}��?	�#����?��)A��?k߰�k�?�$I�$I�?�m۶m��?              �?d!Y�B�?�Mozӛ�?              �?      �?      �?      �?                      �?              �?      �?      �?              �?      �?                      �?      �?      �?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�<�@�0�?d���<�?�'K`�~�?&�i?Y�?��v`��?�%~F��?��8��8�?�q�q�?<<<<<<�?�?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?        t�E]t�?]t�E�?ى�؉��?�؉�؉�?      �?                      �?�������?333333�?�;�;�?�؉�؉�?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?        �������?333333�?�$I�$I�?۶m۶m�?�������?333333�?      �?                      �?d!Y�B�?ӛ���7�?�?�������?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?/�����?	�%��Ю?�������?�?|a���?GX�i��?��I��I�?l�l��?UUUUUU�?UUUUUU�?              �?      �?              �?        w�'�K�?H���@��?              �?�������?�������? �����? �����?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ[س=hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         b                    �?U�ք�?�           ��@              ;       
             �?j�[y۾�?�            y@                     	          ����?�,M���?�            �r@                                   �?\-��p�?C             ]@                                   @M@     ��?             0@                                 �k@�q�q�?             (@        ������������������������       �                      @               	       	          ����?      �?             $@        ������������������������       �                      @        
                          �s@      �?              @                                  �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                  �i@�ڊ�e��?8             Y@       ������������������������       �        "            �N@                                    L@�θ�?            �C@        ������������������������       �                     4@                                  �_@�\��N��?             3@                                 @_@�q�q�?	             .@        ������������������������       �                     @                                   [@�eP*L��?             &@                                  �?r�q��?             @        ������������������������       �                     @                                   @N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               :                   Pe@Hx�i�.�?o             g@               +                    \@x�û��?n             g@        !       &                   �_@x�}b~|�?#            �L@        "       %                    �J@�	j*D�?             *@        #       $       	             @և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        '       (                   @s@`���i��?             F@       ������������������������       �                    �C@        )       *                   �[@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ,       -                    @L@ ���z��?K            �_@        ������������������������       �        !             N@        .       3                    \@0�,���?*            �P@        /       2                   �`@      �?              @        0       1                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        4       5                    c@P����?&            �M@       ������������������������       �        "             K@        6       9                   �a@z�G�z�?             @        7       8                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        <       M                    �L@�JY�8��?C             Y@       =       J       	            �?�θ�?*            @P@       >       ?                    c@���C��?!            �J@       ������������������������       �                     A@        @       A                    �?�����?             3@        ������������������������       �                     @        B       C                     B@և���X�?	             ,@        ������������������������       �                      @        D       I                    �I@�q�q�?             (@       E       H                    �?z�G�z�?             $@       F       G                   �h@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        K       L                    �?      �?	             (@        ������������������������       �                     @        ������������������������       �                     "@        N       a                   `c@<=�,S��?            �A@       O       \                    �?*;L]n�?             >@       P       Q       	          ����?���Q��?             4@        ������������������������       �                     @        R       S                    �?�n_Y�K�?
             *@        ������������������������       �                      @        T       [                    @N@���!pc�?             &@       U       V                    �?      �?             @        ������������������������       �                     �?        W       X                   @_@���Q��?             @        ������������������������       �                      @        Y       Z       	          033�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ]       `                    @M@ףp=
�?             $@        ^       _                   h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        c       t                   �c@���jm��?�            �t@        d       g                    �?��<b���?             G@        e       f                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        h       s                     P@R���Q�?             D@       i       l                    �?�KM�]�?             C@        j       k       	          @33�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        m       n       
             �?�IєX�?             A@       ������������������������       �                     :@        o       r                   �b@      �?              @       p       q                    @J@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        u       �                   �`@d��=���?�            �q@       v       �                    �?Z�ڤ��?}             h@       w       �                    �?����ր�?m            @d@        x       y                   @[@r֛w���?             ?@        ������������������������       �                      @        z       �                   �m@V�a�� �?             =@        {       |                    b@X�Cc�?
             ,@        ������������������������       �                     @        }       ~                    `@�eP*L��?             &@        ������������������������       �                      @               �                   �e@�q�q�?             "@       ������������������������       �                     @        �       �                    �E@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @L@��S�ۿ?
             .@       ������������������������       �                     (@        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?�1����?X            ``@        �       �                   �[@�������?             A@        ������������������������       �                      @        �       �                    �?     ��?             @@       �       �                   d@r�q��?             >@       �       �       	          ��� @�E��ӭ�?             2@       �       �                   �^@     ��?             0@       �       �                   �]@�q�q�?             "@        ������������������������       �                     @        �       �                   @c@      �?             @       �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                      @        �       �                    @`�E���?A            @X@       �       �                   (p@�L��ȕ?>            @W@       ������������������������       �        '             O@        �       �                     L@�g�y��?             ?@       ������������������������       �                     8@        �       �                    �L@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?r֛w���?             ?@        �       �                    @Q@և���X�?             ,@       �       �                    @���Q��?             $@       �       �       	          ����?և���X�?             @        ������������������������       �                      @        �       �                   �p@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     1@        �       �       
             �?���!���?B            �W@        �       �                    �?��P���?            �D@        �       �                    �P@�eP*L��?             &@       �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                   �i@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   Pa@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �R@ףp=
�?             >@       �       �                   8r@ 	��p�?             =@       �       �                   �`@ ��WV�?             :@       ������������������������       �                     7@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@ �h�7W�?&            �J@        ������������������������       �                     7@        �       �                   0c@ףp=
�?             >@        ������������������������       �                      @        �       �                   �c@h�����?             <@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �       	          ����?�q�q�?             @       �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�Bp  ᓔ��?�5�;��?)OD��?=�5��?"8vi�?]��8�r�?�{a���?a����?      �?      �?�������?�������?      �?              �?      �?              �?      �?      �?      �?      �?      �?                      �?      �?                      �?
ףp=
�?��Q��?              �?�؉�؉�?ى�؉��?              �?�5��P�?y�5���?UUUUUU�?UUUUUU�?              �?]t�E�?t�E]t�?�������?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?        @bw�#�?��X���?8��Moz�?-d!Y��?Lg1��t�?�YLg1�?;�;��?vb'vb'�?�$I�$I�?۶m۶m�?              �?      �?                      �?F]t�E�?F]t�E�?              �?�������?�������?              �?      �?        �@ �?�����~�?              �?g��1��?Ez�rv�?      �?      �?      �?      �?      �?                      �?              �?'u_[�?�V'u�?              �?�������?�������?      �?      �?              �?      �?                      �?      �?        )\���(�?�G�z��?ى�؉��?�؉�؉�?\�琚`�?"5�x+��?      �?        Q^Cy��?^Cy�5�?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?                      �?      �?      �?      �?                      �?X|�W|��?�A�A�?�������?""""""�?333333�?�������?      �?        ى�؉��?;�;��?      �?        t�E]t�?F]t�E�?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?              �?Ri�!$��?[-Y����?��Moz��?��,d!�?UUUUUU�?UUUUUU�?      �?                      �?333333�?333333�?(�����?�k(���?      �?      �?              �?      �?        �?�?              �?      �?      �?�������?333333�?      �?                      �?              �?      �?        ���L�?�#(ͦ�?���
���?n����?Ix�5?�?�5?,R�?���{��?�B!��?              �?��{a�?a���{�?%I�$I��?�m۶m��?      �?        t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?        �������?333333�?      �?                      �?�������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        J�eDP�?����?�������?�������?              �?      �?      �?�������?UUUUUU�?�q�q�?r�q��?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?              �?      �?      �?              �?      �?              �?              �?                      �?      �?                      �??��W�?����?��~���?X`��?      �?        ��{���?�B!��?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?���{��?�B!��?۶m۶m�?�$I�$I�?333333�?�������?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?                      �?      �?                      �?      �?        �+���?�٨�l��?�����?������?t�E]t�?]t�E�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?                      �?�������?�������?�{a���?������?;�;��?O��N���?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ��sHM0�?"5�x+��?      �?        �������?�������?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJnխphG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKㅔh��B�8         �       
             �?6������?�           ��@              I                    �?<�'���?
           0{@                                  �g@�1��n�?g            �e@                                  �c@�?�<��?)            @P@                                  �?��a�n`�?'             O@                                  �a@�<ݚ�?             ;@              
                    �?      �?             0@              	       	             �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                      	          `ff�?r�q��?             @                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                    �A@                                  �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               &                   �_@      �?>             [@               %                    �R@�������?             >@              $       	          033�?�>4և��?             <@                                  �M@�n_Y�K�?             *@                                  �I@և���X�?             @        ������������������������       �                     �?                                   �?�q�q�?             @        ������������������������       �                     @                                  8w@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                !                    �P@r�q��?             @       ������������������������       �                     @        "       #                    �Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                      @        '       4       	          833�?���L��?*            �S@        (       -                    @I@      �?             4@        )       ,                    �?ףp=
�?             $@       *       +                   Pn@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        .       /                   �^@���Q��?             $@        ������������������������       �                     @        0       3                    �?؇���X�?             @        1       2                   0d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        5       F       	             @�c�Α�?             M@       6       7                    �G@��[�8��?            �I@        ������������������������       �                     ,@        8       9                     I@V������?            �B@        ������������������������       �                     @        :       A                    �?     ��?             @@        ;       @       	          ����?�q�q�?
             (@       <       ?                   �b@�<ݚ�?             "@        =       >                    _@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        B       C       	          ����?P���Q�?
             4@        ������������������������       �                     $@        D       E       	          ����?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        G       H                     @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        J       K       	          833�?8Ӈ���?�            `p@        ������������������������       �                    �F@        L       Q       	          ����?<J96���?�             k@        M       N       	          hff�?      �?              @        ������������������������       �                      @        O       P                    �L@      �?             @        ������������������������       �                     @        ������������������������       �                     @        R       S                   �Z@�KM�]�?�             j@        ������������������������       �                     @        T                           �?���"F��?�            `i@       U       l                    @L@ ��Ou��?a            �c@       V       e                    �?XB���?4            �U@       W       d       	          ����?�g<a�?-            @S@       X       c                    `@P���Q�?             D@       Y       \                   0g@HP�s��?             9@        Z       [                   �_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ]       b                    �?���7�?             6@        ^       _                    �H@      �?             @        ������������������������       �                      @        `       a                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �        	             .@        ������������������������       �                    �B@        f       k                   �a@ףp=
�?             $@       g       h                    [@z�G�z�?             @       ������������������������       �                     @        i       j                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        m       ~       	          ��� @�θV�?-            @Q@       n       }                    �R@؇���X�?!            �H@       o       p                   �d@      �?              H@        ������������������������       �        
             0@        q       r                   �\@     ��?             @@        ������������������������       �                     @        s       |                    �N@ܷ��?��?             =@        t       u                    @M@�q�q�?             "@        ������������������������       �                     @        v       {                    �?      �?             @       w       z                     N@      �?             @       x       y                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     4@        ������������������������       �                     �?        ������������������������       �                     4@        �       �       	          ����?��E�B��?!            �G@        ������������������������       �                     �?        �       �                   �`@�q��/��?              G@       �       �                   �_@�7��?            �C@        �       �       
             �?      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                    Z@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ?@        �       �                    Z@և���X�?             @        ������������������������       �                      @        �       �                    @G@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?^��˪�?�            �r@        �       �                   �j@����l�?C            @X@        �       �       	          ����?��i#[�?             E@        �       �                    �?�eP*L��?             6@       �       �                    �?X�Cc�?	             ,@        ������������������������       �                      @        �       �                   �b@�q�q�?             (@        ������������������������       �                     @        �       �                   �b@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �d@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   Pe@R���Q�?             4@       �       �                   `b@�KM�]�?             3@       �       �                   @^@�X�<ݺ?             2@        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             (@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �L@x��}�?%            �K@       �       �                   Pb@���H��?             E@       ������������������������       �                     3@        �       �       	          ����?��<b���?             7@       �       �                    `@؇���X�?             5@       �       �                    �?�q�q�?             "@       �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                      @        �       �                   pe@�n_Y�K�?             *@       �       �       	          ����?z�G�z�?             $@        �       �                   hp@�q�q�?             @        ������������������������       �                     �?        �       �                     O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	          033�?���a�\�?            @i@       �       �                     R@��:x�ٳ?{            �h@       �       �                    @ ���J��?z            `h@       �       �                    �?��<b�ƥ?r             g@       �       �                   pa@P�Lt�<�?b             c@       �       �                    @L@@m���?G             ]@       ������������������������       �        >            @Y@        �       �                   �a@��S�ۿ?	             .@        ������������������������       �                     @        �       �                   r@      �?              @       �       �                   0b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pc@�8��8��?             B@       �       �                   �t@�����H�?             ;@       �       �                    �?`2U0*��?             9@        �       �                   �k@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @@        �       �                   �j@�C��2(�?             &@        �       �                    �?�q�q�?             @       �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  ��X�5�?��S�$e�?��A0�?�>���s�?]�����?Q��#��? �����?�����?�c�1Ƹ?�s�9��?�q�q�?9��8���?      �?      �?�������?�������?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?�������?�������?�m۶m��?�$I�$I�?ى�؉��?;�;��?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?      �?        �4H�4H�?��o��o�?      �?      �?�������?�������?�$I�$I�?۶m۶m�?      �?                      �?              �?�������?333333�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?5�rO#,�?�{a���?�?�������?      �?        �g�`�|�?o0E>��?              �?      �?      �?�������?�������?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?ffffff�?�������?      �?        �������?�������?              �?      �?        �$I�$I�?�m۶m��?              �?      �?        ����a�?�*NHɳ�?              �?�h�?ڿ?�p	��?      �?      �?      �?              �?      �?      �?                      �?(�����?�k(���?      �?        ��%f-�?\E;Sz�?�i�i�?.��-���?�{a���?GX�i���?�cj`?���8+�?�������?ffffff�?{�G�z�?q=
ףp�?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?�.�袋�?      �?      �?              �?      �?      �?              �?      �?                      �?              �?              �?�������?�������?�������?�������?              �?      �?      �?      �?                      �?              �?�Q�g���?̵s���?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?        a���{�?��=���?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?      �?                      �?AL� &W�?�l�w6��?      �?        ��Mozӻ?�B����?�A�A�?��[��[�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?�x��S�?��_��?2���$�?��Id��?�<��<��?�a�a�?]t�E�?t�E]t�?%I�$I��?�m۶m��?      �?        �������?�������?      �?        �q�q�?r�q��?      �?                      �?      �?      �?              �?      �?        333333�?333333�?(�����?�k(���?�q�q�?��8��8�?UUUUUU�?�������?      �?                      �?              �?      �?              �?        pX���o�?A��)A�?�0�0�?��y��y�?      �?        ��,d!�?��Moz��?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?ى�؉��?;�;��?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        D�I��A�?��g���?
�����?[�R�֯�?��-��-�?�A�A�?��7��M�?d!Y�B�?���k(�?(�����?�{a��?�{a���?      �?        �������?�?      �?              �?      �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?�q�q�?�q�q�?���Q��?{�G�z�?      �?      �?      �?              �?      �?              �?      �?              �?                      �?      �?              �?        ]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�[�.hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�/         n                    �?��Wޫ��?�           ��@              e                    �?�y#���?�            �x@              @                   �b@(���@��?�            �q@                                  �?      �?�             m@                                  �`@`՟�G��?             ?@                     	          ����?�X�<ݺ?             2@       ������������������������       �                     $@                                  �Z@      �?              @        	       
                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@               '       	          ����?|u#���?{             i@                                  @E@<��¤�?*             Q@                                   �?HP�s��?             9@       ������������������������       �                     2@                                  `Y@����X�?             @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                       
             �?�K��&�?            �E@                                  �k@�t����?             1@        ������������������������       �                      @                                   �?�<ݚ�?             "@                                  @J@      �?              @       ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        !       &                    ]@ȵHPS!�?             :@        "       %                    �?և���X�?             @        #       $                    �N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@        (       9                   @j@�KM�]�?Q            �`@        )       6                    �?ҳ�wY;�?             A@       *       +                    �?�c�Α�?             =@        ������������������������       �                     �?        ,       -                   `_@����X�?             <@        ������������������������       �                     $@        .       /                    `@X�<ݚ�?	             2@        ������������������������       �                     @        0       1                   �W@r�q��?             (@        ������������������������       �                     �?        2       5                    �?�C��2(�?             &@        3       4       	          ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        7       8       	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        :       ;                    `P@��F�D�?;            �X@       ������������������������       �        7            �W@        <       ?                    �?���Q��?             @        =       >                     Q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        A       d       	             @��H�}�?$             I@       B       C                    Z@(���@��?!            �G@        ������������������������       �                      @        D       O                   d@���X�K�?             �F@        E       J       
             �?R���Q�?             4@        F       G                    �?���Q��?             @        ������������������������       �                      @        H       I                    q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        K       N                    �G@��S�ۿ?             .@        L       M                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        P       c                   @c@���Q��?             9@       Q       b                     N@�LQ�1	�?             7@       R       Y                   �d@      �?             4@        S       V       	             �?���Q��?             @       T       U                   m@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        W       X                   0`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Z       a                    k@�r����?             .@        [       `                   �e@�q�q�?             @       \       _       	             �?�q�q�?             @       ]       ^                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        f       k       
             �?���^���?M            �\@       g       h                    y@�a�O�?B            @X@       ������������������������       �        ?            �W@        i       j                   @X@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       m                    @J@b�2�tk�?             2@        ������������������������       �                     @        ������������������������       �                     &@        o       �                    @K@���A��?�            u@       p       �                    �?P���+�?|            �h@       q       �       
             �?�X�<ݺ?m            �f@        r       s                   �Z@���N8�?             E@        ������������������������       �                     @        t       �       	             @:�&���?            �C@       u       |                   �`@�S����?             C@       v       w                    l@�FVQ&�?            �@@        ������������������������       �                     .@        x       y                   �d@�����H�?
             2@        ������������������������       �                     *@        z       {                    @G@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        }       �                    �?z�G�z�?             @        ~                          �g@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        V            @a@        �       �       
             �?�����?             3@       �       �                   �b@�r����?             .@       ������������������������       �        	             *@        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?ڡ�:x��?V            @a@       �       �                   �[@|�i���?0             S@        ������������������������       �                     @        �       �                    �?�1��u�?.            @R@       �       �                    @O@v�2t5�?            �D@       �       �                   �a@�z�G��?             >@        �       �                   �^@�8��8��?             (@        �       �                    Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �`@X�<ݚ�?             2@       �       �                    @L@����X�?             ,@        ������������������������       �                     @        �       �                    �?�C��2(�?             &@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?���!pc�?             &@        ������������������������       �                      @        �       �       	          ����?�����H�?             "@        ������������������������       �                     @        �       �       	          `ff@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �s@     ��?             @@       �       �                    @N@`Jj��?             ?@        ������������������������       �                     0@        �       �                   �`@�r����?
             .@       ������������������������       �                     &@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �^@�n`���?&             O@        ������������������������       �                     $@        �       �                    �?�θ�?!             J@       �       �       	          ��� @Jm_!'1�?             �H@       �       �                     R@�����H�?            �F@       �       �                    �L@Du9iH��?            �E@        �       �                    c@@�0�!��?             1@       �       �                   �^@��S�ۿ?
             .@        ������������������������       �                      @        �       �                   0b@؇���X�?             @        �       �       	          @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     :@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  +^�ɑA�?�P47��?����Ә�?�Ә��?R�٨�l�?W�+���?      �?      �?�1�c��?�s�9��?��8��8�?�q�q�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?��2�?�C��x�?iiiiii�?KKKKKK�?{�G�z�?q=
ףp�?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?��)kʚ�?���)k��?�?<<<<<<�?              �?�q�q�?9��8���?      �?      �?              �?      �?      �?              �?      �?              �?        ��N��N�?�؉�؉�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?              �?        (�����?�k(���?�������?�������?�{a���?5�rO#,�?              �?�$I�$I�?�m۶m��?              �?�q�q�?r�q��?      �?        UUUUUU�?�������?      �?        F]t�E�?]t�E�?      �?      �?              �?      �?                      �?�������?�������?      �?                      �?[�R�֯�?j�J�Z�?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?{�G�z�?
ףp=
�?W�+���?R�٨�l�?              �?l�l��?�'}�'}�?333333�?333333�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�?      �?      �?              �?      �?              �?        333333�?�������?Nozӛ��?d!Y�B�?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �������?�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?              �?                      �?              �?              �?���ϱ?ܯK*��?����? tT����?              �?UUUUUU�?UUUUUU�?      �?                      �?9��8���?�8��8��?      �?                      �?�&�פ�?.���P��?���/M�?�Q7���?��8��8�?�q�q�?�a�a�?��y��y�?              �?�A�A�?�o��o��?(������?^Cy�5�?>����?|���?      �?        �q�q�?�q�q�?      �?        333333�?�������?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?              �?      �?        ^Cy�5�?Q^Cy��?�?�������?              �?      �?              �?        ̵s��?�g��%�?�5��P^�?�5��P�?      �?        �1bĈ�?�s�Ν;�?�ڕ�]��?��+Q��?333333�?ffffff�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?r�q��?�$I�$I�?�m۶m��?      �?        F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?        �������?�������?              �?      �?              �?      �?�B!��?���{��?              �?�?�������?              �?      �?      �?              �?      �?              �?        �9�s��?�c�1��?      �?        ى�؉��?�؉�؉�?����X�?������?�q�q�?�q�q�?qG�w��?w�qGܱ?ZZZZZZ�?�������?�������?�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��=hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�,                            @E@�p9��a�?�           ��@                                   �?@4և���?U            �_@                      
             �?���-T��?(             O@                                   \@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                    M@ܷ��?��?%             M@        ������������������������       �                     :@        	              	          ����?     ��?             @@       
              	             п���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@                      
             �?�eP*L��?             &@                                 �d@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        -             P@               j       	          `ff�?D�n�3��?s            �@              C                    @L@�&���?�            �s@              <                    �?���9yw�?�            �m@                                  �?�NW���?�            �j@        ������������������������       �        1            �S@               +                    �?t�U����?Y            �`@               &                   ``@���!pc�?            �@@                                 �b@�ՙ/�?             5@                                   �?ףp=
�?             $@       ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                !                   j@���|���?	             &@        ������������������������       �                     @        "       %                   �d@և���X�?             @       #       $                   �k@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        '       (                   �n@�8��8��?	             (@       ������������������������       �                     @        )       *                     H@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ,       3                   �]@�L�L��?@            @Y@        -       2                   `\@d}h���?	             ,@       .       /                   �o@�8��8��?             (@       ������������������������       �                     $@        0       1                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        4       ;                    @`��F:u�?7            �U@       5       6                   ``@�D�e���?5            @U@       ������������������������       �                     �I@        7       8                    �?�IєX�?             A@       ������������������������       �                     ;@        9       :                    d@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        =       @                   �b@��}*_��?             ;@       >       ?       
             �?      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        A       B                   0q@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        D       O       
             �?�Q����?0             T@        E       N                    b@���"͏�?            �B@       F       M                   �`@¦	^_�?             ?@       G       H       	          ����?�+$�jP�?             ;@       ������������������������       �        	             1@        I       L                   �b@      �?             $@       J       K                   `b@����X�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        P       Y                   �b@��V#�?            �E@        Q       T                    �L@�q�q�?             8@        R       S                   @]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        U       X                    �?ףp=
�?             4@        V       W                     Q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@        Z       _                   �c@�\��N��?             3@        [       \                    �N@z�G�z�?             @        ������������������������       �                      @        ]       ^                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        `       e                   �q@X�Cc�?             ,@       a       d                   Pd@؇���X�?             @        b       c                    @M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        f       g                   d@և���X�?             @        ������������������������       �                      @        h       i                   `u@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        k       �       	          033�?BSf���?�            r@        l       }                    �?j���� �?:            @U@        m       n                    �G@"pc�
�?            �@@        ������������������������       �                      @        o       p                    @H@�+e�X�?             9@        ������������������������       �                      @        q       |                    �?�㙢�c�?             7@       r       {                    �?������?             1@       s       v                   `]@����X�?             ,@        t       u       	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        w       z                    �?ףp=
�?	             $@        x       y                   �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ~       �                    �?8�Z$���?!             J@              �                    �K@�����?             E@        ������������������������       �                     6@        �       �                   �_@z�G�z�?             4@       �       �                   �\@@4և���?	             ,@        ������������������������       �                     �?        ������������������������       �                     *@        �       �                   Pa@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?���Q��?             $@        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                   `Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �a@L紂P�?r            �i@       �       �       	          pff�?hڛ�ʚ�?V            �b@        �       �                    ]@@4և���?             <@        ������������������������       �                      @        ������������������������       �                     :@        �       �                    \@��7�K¨?E            @^@        �       �                    �?��p\�?            �D@       �       �                   �_@ 7���B�?             ;@        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �                   �c@؇���X�?             ,@        ������������������������       �                     $@        �       �                   �[@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        -             T@        �       �                   �`@<|ۤ$�?            �K@        �       �                   �m@�ՙ/�?             5@       �       �                    �?     ��?             0@       ������������������������       �                     $@        �       �                   `e@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �F@�t����?             A@        ������������������������       �                     @        �       �                    c@��a�n`�?             ?@        �       �                    @�IєX�?             1@       ������������������������       �                     0@        ������������������������       �                     �?        �       �       	             @և���X�?             ,@       �       �                     K@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  !0u(���?�g��29�?�$I�$I�?n۶m۶�?�RJ)���?[k���Z�?      �?      �?              �?      �?        a���{�?��=���?              �?      �?      �?�a�a�?��y��y�?      �?                      �?]t�E�?t�E]t�?�$I�$I�?۶m۶m�?              �?      �?              �?                      �?���k(�?��k(��?Y/�y�?���B�?��Y��?���s��?萚`���?�x+�R�?      �?        ���-�?g��1��?F]t�E�?t�E]t�?�<��<��?�a�a�?�������?�������?      �?              �?      �?      �?                      �?F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?)0��<��?�~�X��?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�u�7[��?Ȥx�L��???????�?�?      �?        �?�?      �?        �m۶m��?�$I�$I�?      �?                      �?              �?B{	�%��?_B{	�%�?      �?      �?              �?      �?        /�袋.�?F]t�E�?      �?                      �?ffffff�?�������?*�Y7�"�?v�)�Y7�?�RJ)���?��Zk���?B{	�%��?/�����?              �?      �?      �?�$I�$I�?�m۶m��?      �?                      �?      �?              �?                      �?eMYS֔�?6eMYS��?UUUUUU�?�������?      �?      �?      �?                      �?�������?�������?      �?      �?              �?      �?              �?        y�5���?�5��P�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?%I�$I��?�m۶m��?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?        `�}2��?躍`3�?ZZZZZZ�?�������?/�袋.�?F]t�E�?      �?        R���Q�?���Q��?              �?�7��Mo�?d!Y�B�?xxxxxx�?�?�m۶m��?�$I�$I�?      �?      �?      �?                      �?�������?�������?      �?      �?      �?                      �?      �?              �?              �?        ;�;��?;�;��?�a�a�?=��<���?              �?�������?�������?�$I�$I�?n۶m۶�?      �?                      �?      �?      �?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?7`��c.�?�y����?�$I�$I�?n۶m۶�?      �?                      �?���!pc�?�0�~�4�?��+Q��?�]�ڕ��?h/�����?	�%����?�$I�$I�?۶m۶m�?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?��7�}��?��)A��?�<��<��?�a�a�?      �?      �?      �?              �?      �?      �?                      �?              �?�������?�������?      �?        �s�9��?�c�1��?�?�?              �?      �?        ۶m۶m�?�$I�$I�?333333�?�������?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��(hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKӅ�h��B�4         x                    �?������?�           ��@              q                   �c@�q��?�             x@              h                    �?���6�?�            �u@              +                    �?b�sG�?�             o@                      
             �?"Mw����?2            @U@                                  �?RB)��.�?            �E@                                 �p@z�G�z�?             D@                                  �?�t����?             A@        	                          �m@և���X�?             @       
                          �R@���Q��?             @        ������������������������       �                     �?                      	          ����?      �?             @        ������������������������       �                     �?                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@                                   �?      �?             @                                  @a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  r@      �?             @        ������������������������       �                     �?                                  �u@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               *                   �c@r�q��?             E@               )                    �G@      �?             D@        !       "                   `]@�q�q�?             .@        ������������������������       �                     @        #       $                   @`@�eP*L��?             &@        ������������������������       �                     @        %       &                   �a@      �?              @       ������������������������       �                     @        '       (                   @`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     9@        ������������������������       �                      @        ,       C       	          ����?�i����?m            �d@        -       0                    �?�Gi����?            �B@        .       /                   �n@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        1       8                   @a@X�Cc�?             <@        2       3                    �?�8��8��?
             (@       ������������������������       �                     "@        4       5                   �^@�q�q�?             @        ������������������������       �                     �?        6       7                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        9       B                   �c@     ��?
             0@       :       ?                   �Z@�	j*D�?             *@        ;       <                   �[@���Q��?             @        ������������������������       �                      @        =       >       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        @       A                   �a@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        D       O       	          ����?R�xE��?V            �_@        E       J                    �?d}h���?             <@       F       I                    �?���N8�?             5@        G       H                   ``@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        K       N                    [@����X�?             @        L       M                    @K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        P       Q                    �?�FVQ&�?D            �X@        ������������������������       �                     *@        R       g                    @N@Du9iH��??            �U@       S       `                   `j@ȵHPS!�?)             J@        T       U       	          033�?����X�?             ,@        ������������������������       �                      @        V       W                    \@�q�q�?             (@        ������������������������       �                      @        X       _                    @M@z�G�z�?	             $@       Y       Z                    _@�����H�?             "@        ������������������������       �                     @        [       \                    �C@z�G�z�?             @        ������������������������       �                     @        ]       ^                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        a       b                     M@�}�+r��?             C@       ������������������������       �                     @@        c       f                    �?�q�q�?             @       d       e                   �`@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     A@        i       j       
             �?�7��d��?B             Y@       ������������������������       �        5            �S@        k       l                    �I@�q�q�?             5@        ������������������������       �                     @        m       p                    �?      �?	             0@        n       o                   �`@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        r       w       	          pff�?����X�?            �A@       s       v                    �M@r٣����?            �@@       t       u                    �? ��WV�?             :@       ������������������������       �                     9@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        y       �                    �?
�:7���?�            �u@       z       �                   `R@2�����?�            @r@        {       |                   �Z@     ��?	             0@        ������������������������       �                     @        }       �                    `@�q�q�?             (@       ~       �                    �?      �?              @              �                   �a@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @r�q��?�            @q@       �       �       
             �?L.��:��?�            @o@        �       �                    �?�xGZ���?'            �Q@        �       �                    c@�θ�?             :@       �       �                   �Z@r�q��?             8@        ������������������������       �                      @        �       �       	          ����?�C��2(�?
             6@        ������������������������       �                     *@        �       �                   @q@�<ݚ�?             "@       ������������������������       �                     @        �       �       	          `ff�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @L@8�A�0��?             F@       �       �                    �I@���Q��?             9@       �       �                     G@j���� �?             1@       �       �                   o@�z�G��?             $@       ������������������������       �                     @        �       �                   �e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	          `ff�?�S����?             3@       �       �       	          ����?�z�G��?             $@       �       �                   �a@؇���X�?             @        ������������������������       �                     @        �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                     L@����?�?t            �f@       ������������������������       �        e             c@        �       �                    �?PN��T'�?             ;@       �       �                    �?��2(&�?             6@        �       �                   �_@      �?              @        ������������������������       �                      @        �       �                    �L@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        �       �                   @r@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?�n_Y�K�?             :@       �       �                    �?���y4F�?             3@       �       �                   �p@�q�q�?	             (@       �       �       	          ����?z�G�z�?             $@       ������������������������       �                     @        �       �                   �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@8^s]e�?'             M@       �       �                    �?t/*�?            �G@        �       �                   �t@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   j@���H��?             E@        ������������������������       �                     6@        �       �       	          `ff�?      �?             4@       �       �       
             �?      �?             $@       �       �       	          ����?      �?              @        ������������������������       �                     @        �       �                   �^@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �t�b�      h�h)h,K ��h.��R�(KK�KK��hb�B0  �sF�v
�?�\��z�?�����*�?�����j�?`�tՁ��?�ע���?��g3�?�?�L� ��?�������?�������?���)k��?S֔5eM�?ffffff�?ffffff�?�?<<<<<<�?�$I�$I�?۶m۶m�?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?      �?      �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?        t�E]t�?]t�E�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�+Q��?��+Q��?#�u�)��?o0E>��?r�q��?�q�q�?      �?                      �?�m۶m��?%I�$I��?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?vb'vb'�?;�;��?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?��`0�?>������?۶m۶m�?I�$I�$�?�a�a�?��y��y�?UUUUUU�?�������?      �?                      �?              �?�m۶m��?�$I�$I�?      �?      �?              �?      �?              �?        |���?>����?              �?w�qGܱ?qG�w��?�؉�؉�?��N��N�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?�q�q�?�q�q�?              �?�������?�������?              �?      �?      �?              �?      �?              �?        (�����?�5��P�?              �?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?              �?�Q���?��(\���?              �?UUUUUU�?UUUUUU�?      �?              �?      �?�$I�$I�?�m۶m��?              �?      �?                      �?�m۶m��?�$I�$I�?>���>�?|���?O��N���?;�;��?      �?                      �?              �?              �?��M�!�?���d���?8p���?ȏ?~��?      �?      �?              �?�������?�������?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?              �?      �?        �������?UUUUUU�?1�Zd�?;�O��n�?�_�_�?�A�A�?ى�؉��?�؉�؉�?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?        9��8���?�q�q�?      �?              �?      �?              �?      �?                      �?/�袋.�?颋.���?333333�?�������?ZZZZZZ�?�������?ffffff�?333333�?      �?              �?      �?              �?      �?                      �?      �?        ^Cy�5�?(������?333333�?ffffff�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?��I��I�?l�l��?      �?        &���^B�?h/�����?��.���?t�E]t�?      �?      �?              �?�������?UUUUUU�?              �?      �?              �?        �������?�������?      �?                      �?;�;��?ى�؉��?6��P^C�?(������?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?	�=����?|a���?W�+���?�;����?333333�?�������?      �?                      �?��y��y�?�0�0�?              �?      �?      �?      �?      �?      �?      �?              �?333333�?�������?      �?                      �?      �?                      �?]t�E�?F]t�E�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���~hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�*         d       
             �?T8���?�           ��@                                  �?�K�x�v�?           �y@                                  �b@r�q��?,             R@                                  �?�D��?            �H@               
                   �\@�q�����?             9@               	                   �q@�<ݚ�?             "@                     
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                      
             �?      �?             0@        ������������������������       �                     @                                   @�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @                                  `a@ �q�q�?             8@       ������������������������       �                     0@                                    K@      �?              @                                  �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?�LQ�1	�?             7@                                  @C@�C��2(�?             6@        ������������������������       �                     �?                                  �b@���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?        ������������������������       �                     �?               +                   �f@���4��?�            0u@                                    �?     ��?K             `@       ������������������������       �        6            �W@        !       *                    �?�IєX�?             A@        "       )                   �`@�r����?	             .@       #       (                    �?����X�?             @       $       '       	          `ff�?      �?             @       %       &                   �X@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@        ,       A                    �?ė���w�?�            `j@        -       2       	          833�?�w�"w��?.             S@        .       1                    a@�nkK�?             7@        /       0                    �E@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     &@        3       4                    ]@䯦s#�?             �J@        ������������������������       �                     @        5       :                   �a@�[�IJ�?            �G@        6       9       	          033�?ףp=
�?             4@        7       8                   8w@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@        ;       @                   @b@�q�q�?             ;@       <       ?                   �d@�û��|�?             7@       =       >                   hp@      �?	             0@       ������������������������       �                     ,@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        B       a                    @Tۢ��(�?^            �`@       C       H                    @G@����?\            @`@        D       G                    �?�θ�?	             *@       E       F                    �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                      @        I       J                   @Z@@\�*��?S            @]@        ������������������������       �                     �?        K       X       	          ����?XB���?R             ]@        L       O                   �\@     ��?             @@        M       N                     N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        P       S                   @X@ 	��p�?             =@        Q       R                   0j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        T       U                    @N@ ��WV�?             :@       ������������������������       �                     .@        V       W                   �`@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        Y       Z                    �? ��N8�?9             U@       ������������������������       �        ,             P@        [       `                    �?P���Q�?             4@       \       _                   ``@�C��2(�?             &@        ]       ^                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        b       c                    �I@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        e       r                   Pc@BK"(<\�?�            0t@        f       m       	            �?�������?             >@        g       h                   �\@      �?              @        ������������������������       �                     �?        i       l                    �?؇���X�?             @        j       k                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        n       q                   @^@���7�?             6@        o       p                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        s       �                    �?�y��>�?�            Pr@       t       �                    �?@9G��?�            �n@        u       �                   �q@ȵHPS!�?$             J@       v       �       	          ����?���}<S�?              G@       w       �                   �l@������?            �D@       x                          �l@PN��T'�?             ;@       y       ~       	          ����?HP�s��?             9@       z       }                   �e@ �q�q�?             8@        {       |                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �D@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�X-:oȤ?v             h@        ������������������������       �        /            �U@        �       �                   �t@PԱ�l�?G            �Z@       �       �                    �?P�c0"�?F            @Z@        �       �                   �b@@4և���?             ,@       ������������������������       �        
             &@        �       �                   `c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    _@@��,B�?:            �V@        �       �       	            �?�Ń��̧?             E@       ������������������������       �                    �A@        �       �       	          pff�?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        #            �H@        ������������������������       �                      @        �       �       	          pff�?     ��?             H@       �       �                    �?8^s]e�?             =@        ������������������������       �                      @        �       �                    `@և���X�?             5@        �       �                   `_@�<ݚ�?             "@       �       �                    �O@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    h@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �       	          033�?�}�+r��?
             3@        �       �                   q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�
  6n����?�� ���?;s�����?1������?UUUUUU�?UUUUUU�??4և���?������?���Q��?�p=
ף�?�q�q�?9��8���?      �?      �?      �?                      �?      �?              �?      �?              �?ى�؉��?�؉�؉�?      �?                      �?UUUUUU�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?��Moz��?Y�B��?]t�E�?F]t�E�?              �?��y��y�?�a�a�?      �?                      �?              �?�Κ�?#��+b��?      �?     ��?              �?�?�?�?�������?�$I�$I�?�m۶m��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?              �?H��i�?.~��%�?��k(��?���k(�?d!Y�B�?�Mozӛ�?UUUUUU�?UUUUUU�?      �?                      �?              �?�V�9�&�?�����?              �?m�w6�;�?���
b�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?8��Moz�?��,d!�?      �?      �?      �?                      �?              �?      �?        �M1j�۴?Hֹ�d�? �����?~�~��?�؉�؉�?ى�؉��?F]t�E�?]t�E�?              �?      �?              �?        ^�^�?���?      �?        �{a���?GX�i���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �{a���?������?UUUUUU�?UUUUUU�?      �?                      �?;�;��?O��N���?              �?F]t�E�?]t�E�?              �?      �?        �a�a�?�y��y��?              �?�������?ffffff�?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?              �?333333�?�������?              �?      �?        �6)D�?3@%[���?�������?�������?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        F]t�E�?�.�袋�?�$I�$I�?۶m۶m�?              �?      �?                      �?������?���E�)�?������?9/���?��N��N�?�؉�؉�?ӛ���7�?d!Y�B�?�|����?������?&���^B�?h/�����?q=
ףp�?{�G�z�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �_��7V�?��H	9�?      �?        �N]����?�+J�#�??�c?�c�?8�8��?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        `��_���?h�h��?��<��<�?�a�a�?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?                      �?      �?      �?|a���?	�=����?      �?        �$I�$I�?۶m۶m�?�q�q�?9��8���?�������?333333�?      �?                      �?              �?�������?UUUUUU�?              �?      �?        (�����?�5��P�?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJCLUhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKÅ�h��B�0         �                    �?0����?�           ��@              u                    �?눘ķ�?           �|@              f       	          033�?6�v[X�?�             w@                                 �c@�?6ˠ��?�             t@                                   �N@\�Uo��?             C@                     	             �?      �?             >@                     	          ����?���Q��?             9@              	       
             �?�eP*L��?             6@        ������������������������       �                     "@        
                           �?$�q-�?             *@       ������������������������       �                      @                      	            �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @               5                    �?v^|�_�?�            �q@               4                    �?�.�+��?4            �U@              !       
             �?�w�r��?-            @S@                                   �?���>4��?             <@                                   @O@"pc�
�?             &@       ������������������������       �                      @                                   `P@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                   `@������?             1@        ������������������������       �                     $@                                   �`@և���X�?             @                     	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        "       1       	          833�?���c�H�?            �H@       #       (                    �I@�������?             F@       $       '                    �D@@4և���?             <@        %       &                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     4@        )       0                    `@     ��?             0@       *       /                   �c@      �?             (@       +       ,                   �l@ףp=
�?             $@       ������������������������       �                     @        -       .                   �p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        2       3                    o@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        6       7                   `X@LT���Y�?v            �h@        ������������������������       �                      @        8       ]                   �b@���Ls�?u            `h@       9       N       
             �? 
��р�?h             e@        :       ;                   �j@z�G�z�?            �A@        ������������������������       �                     (@        <       C       	          ����?8����?             7@        =       @                    �?      �?             $@        >       ?                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        A       B                   Pc@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        D       E       	          ����?8�Z$���?             *@        ������������������������       �                     @        F       G       	          ����?      �?              @        ������������������������       �                     �?        H       M                   @c@؇���X�?             @        I       J                    _@�q�q�?             @        ������������������������       �                     �?        K       L       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        O       P                   �^@��J��i�?P            �`@        ������������������������       �        %             P@        Q       R                     L@hA� �?+            �Q@       ������������������������       �        $            �L@        S       T                     M@�θ�?             *@        ������������������������       �                     �?        U       V                    �?r�q��?             (@        ������������������������       �                     @        W       X                    a@      �?              @        ������������������������       �                     �?        Y       Z                    �?؇���X�?             @        ������������������������       �                     @        [       \                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                    �H@�	j*D�?             :@        ������������������������       �                     @        `       a                    �?��<b���?             7@        ������������������������       �                     $@        b       c                    �?�n_Y�K�?             *@        ������������������������       �                     @        d       e                   @_@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        g       p       
             �?���j��?             G@       h       k                    �G@4?,R��?             B@        i       j                   0a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        l       m                    @      �?             @@       ������������������������       �                     8@        n       o                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        q       r                   `U@z�G�z�?             $@        ������������������������       �                     �?        s       t                   �d@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        v       {       
             �?Z��:���?7            �V@       w       z       
             �?�h����?"             L@        x       y                   @_@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     G@        |       �       	          ����?��R[s�?            �A@       }       ~                   �`@$�q-�?             :@       ������������������������       �                     (@               �                   @b@؇���X�?             ,@        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @b@�<ݚ�?             "@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?H%u��?�            0q@        �       �                    �?�D��??            �X@       �       �       
             �?������?4            @U@       �       �                    �?��IF�E�?(            �P@       �       �                   �l@���7�?             F@        ������������������������       �                     9@        �       �       	          ����?�KM�]�?             3@       �       �                   �b@�<ݚ�?             "@       �       �       	          433�?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �       	             �?�GN�z�?             6@        ������������������������       �                     $@        �       �                    @K@�q�q�?             (@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                    �?����X�?             @        ������������������������       �                      @        �       �                    �N@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	             �?�����?             3@       �       �                   �Z@؇���X�?	             ,@        ������������������������       �                     �?        �       �                    h@$�q-�?             *@        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   @`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `P@��
ц��?             *@       �       �                   �`@���|���?
             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   Pj@���r�?v             f@        ������������������������       �        '             P@        �       �                   �j@ (��?O            @\@        ������������������������       �                      @        �       �                    �?�ܗ1�?N            �[@       �       �                   Xq@�zvܰ?=             V@       �       �                   q@ "��u�?"             I@       �       �       	             �?�Ń��̧?             E@        �       �                    @I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �C@        �       �                   0`@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     C@        �       �                    �R@���}<S�?             7@       ������������������������       �                     5@        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  ���^L�?���Y�?u�u��?k�k��?��Moz��?�,d!Y�?��p��?�l<�?�?�5��P^�?6��P^C�?      �?      �?333333�?�������?t�E]t�?]t�E�?              �?�؉�؉�?;�;��?      �?        �������?�������?      �?                      �?      �?                      �?      �?        $Zas ��?p�z2~��?�f��o�?�2)^ �?{����1�?
qV~B��?n۶m۶�?I�$I�$�?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?xxxxxx�?              �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?              �?        4և����?/�����?t�E]t�?/�袋.�?n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?              �?      �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?333333�?�������?      �?                      �?      �?        ��*S��?J�f��?              �?�����?z�z��?	j*D�?�n_Y�K�?�������?�������?      �?        d!Y�B�?8��Moz�?      �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ;�;��?;�;��?      �?              �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        �[�՘H�?���@��?      �?        ���?_�_�?      �?        ى�؉��?�؉�؉�?              �?�������?UUUUUU�?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        vb'vb'�?;�;��?              �?��,d!�?��Moz��?      �?        ;�;��?ى�؉��?      �?        �$I�$I�?�m۶m��?      �?                      �?!Y�B�?ozӛ���?r�q��?�8��8��?      �?      �?              �?      �?              �?      �?              �?      �?      �?      �?                      �?�������?�������?              �?�q�q�?�q�q�?      �?                      �?TFeTFe�?�\��\��?۶m۶m�?�$I�$I�?333333�?ffffff�?              �?      �?                      �?X|�W|��?PuPu�?�؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?        �m۶m��?�$I�$I�?              �?      �?        �q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?        ���Q��?)\���(�??4և���?������?�?xxxxxx�?'�l��&�?�l��&��?F]t�E�?�.�袋�?              �?(�����?�k(���?�q�q�?9��8���?      �?      �?              �?      �?              �?                      �?]t�E�?�袋.��?              �?�������?�������?              �?      �?      �?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?                      �?              �?Q^Cy��?^Cy�5�?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?                      �?�؉�؉�?�;�;�?F]t�E�?]t�E]�?              �?      �?              �?        �^o�?�?�
���?              �?x�!���?H���?      �?        q��$�?�蕱���?t�E]t�?颋.���?���Q��?�G�z�?�a�a�?��<��<�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?                      �?d!Y�B�?ӛ���7�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKۅ�h��B�6         Z                   �`@
���P��?�           ��@               G       
             �?���{��?�            �s@                                  �?d��cό�?�             o@                                   @�����?             3@                                 �v@������?             1@                                 @[@����X�?             ,@        ������������������������       �                     @                                  �n@      �?              @        	       
                    �Q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                      	          ���@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @               F                   �z@t��%�?�            �l@              3                    �?��^ҺR�?�            �l@              (                   ``@P�9�׸?s             f@                                   @O@pH����?.            �P@                                 �[@�h����?&             L@                                   �K@      �?             0@       ������������������������       �                     "@                                  �^@����X�?             @       ������������������������       �                     @        ������������������������       �                      @                                  �X@�(\����?             D@                                  0j@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �A@                '                   `]@���|���?             &@       !       &                    �?�<ݚ�?             "@       "       #                    _@�q�q�?             @        ������������������������       �                      @        $       %                   �Z@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        )       2                   �l@����q�?E            @[@       *       1                   pl@Pa�	�?(            �P@       +       0                    �D@ ����?'            @P@        ,       -                    _@�q�q�?             @        ������������������������       �                     �?        .       /                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        $             O@        ������������������������       �                     �?        ������������������������       �                    �E@        4       A                   �c@�T`�[k�?            �J@       5       @                   �s@�p ��?            �D@       6       9                    �?�˹�m��?             C@       7       8                   �X@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        :       ;       
             �?�t����?	             1@        ������������������������       �                     @        <       ?                   `^@"pc�
�?             &@        =       >       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        B       C       	          ����?      �?             (@        ������������������������       �                     @        D       E                   �d@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        H       Q                    �?���e��?*            �P@       I       L                   @c@r�q��?             E@        J       K       	          433�?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        M       N                    @Pa�	�?            �@@       ������������������������       �                     >@        O       P       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        R       Y                   �c@      �?             8@       S       X                    �?ҳ�wY;�?             1@       T       W                     O@d}h���?	             ,@       U       V                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        [       �       
             �?����T�?�            0z@        \       {                   �_@b�/#w�?i            �d@        ]       f                    �?     ��?'             P@        ^       e                   `]@��2(&�?             6@       _       `                   �k@z�G�z�?             .@        ������������������������       �                     @        a       d       	          ����?      �?              @       b       c                    �D@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        g       l                   �a@����X�?             E@        h       k                    ]@      �?              @        i       j                   j@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        m       n                    Z@H�V�e��?             A@        ������������������������       �                     �?        o       x       	          033�?"pc�
�?            �@@       p       q                   �]@ 7���B�?             ;@        ������������������������       �                     $@        r       s       	          ����?�IєX�?             1@       ������������������������       �                     ,@        t       w                    �?�q�q�?             @       u       v                    o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        y       z                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        |       �                    �?�ެD��?B            �Y@        }       �                   �a@      �?             @@       ~                           �J@�q�q�?             8@       ������������������������       �                     .@        �       �       	          @33�?�����H�?             "@       ������������������������       �                     @        �       �                    a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     E@�ӖF2��?/            �Q@        �       �                    �C@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�? Da�?,            �O@       �       �                    �L@�?�|�?            �B@        �       �                   �h@�IєX�?             1@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �                     4@        �       �                    d@R�}e�.�?             :@       �       �                     O@"pc�
�?             6@       �       �                   �r@�t����?             1@       �       �                    �?      �?             0@        �       �                    @K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     �?        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �L@r�q��?�            �o@       �       �                    �?<2r�Y�?t             h@       �       �                    @L@���#�İ?i             f@       �       �                    �?0)�ci��?f            �e@        �       �       	            �?�����H�?             B@       �       �                   `\@(;L]n�?             >@        �       �                   �[@ףp=
�?             $@       ������������������������       �                      @        �       �                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    �G@      �?             @       �       �       	          hff�?      �?             @        ������������������������       �                      @        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �       	             @�Ŗ�Pw�?Q            @a@       ������������������������       �        P             a@        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?     ��?             0@       �       �       	          ����?      �?             (@       �       �                   �Y@      �?             @        ������������������������       �                      @        �       �                    @K@      �?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                     P@����*��?!            �M@       �       �                    `@�D����?             E@        �       �       	          ����?�q�q�?             (@        ������������������������       �                     @        �       �                    a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �M@�z�G��?             >@        �       �       	          ����?�	j*D�?             *@        ������������������������       �                     @        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     1@        �       �                    �?�t����?             1@       ������������������������       �        	             ,@        �       �                     R@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  փmM���?>IY�8�?��	��	�?ُ�؏��?�����ɼ?�A���f�?^Cy�5�?Q^Cy��?�?xxxxxx�?�$I�$I�?�m۶m��?              �?      �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?              �?      �?        �q�.�|�?�(�j��?����y�?��G���?/�袋.�?]t�E]�?z�rv��?�1���?۶m۶m�?�$I�$I�?      �?      �?              �?�$I�$I�?�m۶m��?              �?      �?        �������?333333�?�������?�������?      �?                      �?              �?F]t�E�?]t�E]�?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?        �,�M�ɒ?���%�i�?|���?|���? �����? �����?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?                      �?"5�x+��?���!5��?��+Q��?Q��+Q�?^Cy�5�?��P^Cy�?�a�a�?��y��y�?      �?                      �?�?<<<<<<�?              �?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?        �>���?>���>�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?|���?|���?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�������?�������?۶m۶m�?I�$I�$�?      �?      �?              �?      �?                      �?      �?                      �?���ڞ�?���J��?E���w��?^�/7Ā�?     ��?      �?t�E]t�?��.���?�������?�������?              �?      �?      �?333333�?�������?              �?      �?                      �?              �?�m۶m��?�$I�$I�?      �?      �?333333�?�������?      �?                      �?              �?iiiiii�?ZZZZZZ�?              �?/�袋.�?F]t�E�?	�%����?h/�����?      �?        �?�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        UUUUUU�?�������?              �?      �?        ��`����?��O ���?      �?      �?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�z2~���?Zas �
�?      �?      �?              �?      �?        AA�?�������?к����?*�Y7�"�?�?�?      �?      �?      �?                      �?              �?              �?�;�;�?'vb'vb�?F]t�E�?/�袋.�?�?<<<<<<�?      �?      �?      �?      �?      �?                      �?              �?      �?        �������?333333�?              �?      �?              �?      �?      �?                      �?�������?UUUUUU�?"fs�P��?��d�x�?��N��?'u_[�?�I���?��֡�l�?�q�q�?�q�q�?�������?�?�������?�������?      �?              �?      �?      �?                      �?      �?              �?      �?      �?      �?              �?      �?      �?              �?      �?              �?        ��?���?ہ�v`�}?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?      �?      �?      �?      �?              �?      �?      �?      �?      �?              �?      �?              �?                      �?      �?        'u_[�?�A�I�?z��y���?�0�0�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?333333�?ffffff�?vb'vb'�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?<<<<<<�?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ"�a,hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@>         z       	          ����?4�5����?�           ��@              G                    �K@t$*�J�?�            �w@              8                    �?��ga�=�?�            �p@              	                   @[@�P��G7�?�            @m@                                  @W@�8��8��?             (@                                  �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        
       -                    �?b�����?�            �k@                                  �?�G�V�e�?~            �i@                                  �Q@��?^�k�?*            �Q@        ������������������������       �                      @        ������������������������       �        )             Q@                                  �c@X�@��l�?T            �`@                                  c@�n_Y�K�?             *@                                  �?r�q��?             @                                  P@      �?             @                      	          �����      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                    �?d�.����?L            @^@                      
             �?���Q��?            �A@        ������������������������       �                     *@                                  �[@���7�?             6@                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        !       *                    @��+��<�?6            �U@       "       )       	          ����?�Ń��̧?4             U@       #       (                   �a@��'�`�?3            �T@        $       %                   `a@���N8�?             5@       ������������������������       �                     3@        &       '                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        &             O@        ������������������������       �                     �?        +       ,                    q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        .       /                   �g@X�<ݚ�?             2@        ������������������������       �                     @        0       1                     C@r�q��?	             (@        ������������������������       �                     �?        2       3                   �n@�C��2(�?             &@       ������������������������       �                     @        4       5                    ^@      �?             @        ������������������������       �                      @        6       7                    p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        9       :                   �U@j���� �?             A@        ������������������������       �                     $@        ;       @                    �?r�q��?             8@       <       =                    �?�IєX�?             1@       ������������������������       �        
             .@        >       ?                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        A       B                   @^@և���X�?             @        ������������������������       �                      @        C       D                    �?���Q��?             @        ������������������������       �                     �?        E       F       	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        H       s                    �?��7Y��?N            �[@       I       ^       
             �?|��?���?:            @T@        J       [                   �d@�<ݚ�?             B@       K       X       	          ����?     ��?             @@       L       U                   �p@$�q-�?             :@       M       T                   �X@ �q�q�?             8@        N       S                    �?      �?              @       O       P                    �?r�q��?             @        ������������������������       �                     @        Q       R                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        V       W                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                     O@      �?             @        ������������������������       �                     @        ������������������������       �                     @        \       ]                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        _       n                    �?f.i��n�?            �F@       `       m                    �?��
ц��?             :@       a       l                   @a@���Q��?             4@       b       k                    `P@և���X�?             ,@       c       j                    �?�q�q�?	             (@       d       e                   �k@z�G�z�?             $@       ������������������������       �                     @        f       i       	          ����?�q�q�?             @       g       h                   �s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        o       p       	            �?�KM�]�?             3@       ������������������������       �                     ,@        q       r                    q@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        t       u       
             �?�������?             >@       ������������������������       �                     2@        v       y                   @b@�q�q�?             (@       w       x                    Z@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        {       �                    �?ܫV�L%�?�            0v@        |       �                    �?     8�?%             P@       }       �                    �?:ɨ��?            �@@        ~       �                   pp@      �?	             ,@              �                    �E@�z�G��?             $@        ������������������������       �                     �?        �       �       
             �?�<ݚ�?             "@        ������������������������       �                     �?        �       �       
             �?      �?              @       �       �                   `g@z�G�z�?             @        ������������������������       �                      @        �       �                   @_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   `^@�S����?
             3@        �       �                   �`@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        �       �                   �c@��� ��?             ?@       �       �                    �?h�����?             <@        ������������������������       �                     "@        �       �                    �K@�}�+r��?             3@       ������������������������       �                     (@        �       �                    q@؇���X�?             @       ������������������������       �                     @        �       �                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �v@�Ι����?�            0r@       �       �       
             �?P�I;l�?�            �q@       �       �                    f@L���?�            @n@       �       �                    �?\ ���?�            �m@        �       �       	          ����?���-T��?*             O@        �       �                     L@X�Cc�?             ,@        �       �                   �[@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     E@�8��8��?             H@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   d@���.�6�?             G@       �       �       	          `ff�? �#�Ѵ�?            �E@        �       �                   �b@؇���X�?
             ,@       �       �                     M@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     =@        �       �       	          `ff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �R@(��z�(�?p            �e@       �       �                    �?���1j	�?n            �e@       �       �                   @_@���N8�?^            `b@        �       �                   �_@ȵHPS!�?             :@       �       �                   �^@     ��?             0@       �       �                    �K@�8��8��?	             (@       ������������������������       �                      @        �       �       
             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ���@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        �       �                   pa@Xsj�]�?J            @^@        ������������������������       �                     C@        �       �                   �e@��`qM|�?/            �T@        �       �                   pb@�r����?	             .@        ������������������������       �                     @        �       �                   `U@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                    q@г�wY;�?&             Q@       ������������������������       �                     E@        �       �                   Xq@$�q-�?             :@        ������������������������       �                      @        ������������������������       �                     8@        �       �                    �?H%u��?             9@        ������������������������       �                     �?        �       �       	             �?�8��8��?             8@        �       �                   �`@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             0@        �       �                   �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�4F����?            �D@        �       �                    @F@�\��N��?             3@        ������������������������       �                      @        �       �                    �J@��.k���?             1@        ������������������������       �                     @        �       �                    �?�n_Y�K�?	             *@        ������������������������       �                     �?        �       �       	          ���@�q�q�?             (@       �       �                    d@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �^@��2(&�?             6@        �       �                    �?���Q��?             @       �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�IєX�?             1@       ������������������������       �        	             .@        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �a@      �?              @       �       �                   ``@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �t�b�
     h�h)h,K ��h.��R�(KK�KK��hb�B�   Np	�?���Gw{�?�A-'r�?��|���?��[���?�1���?Z��Y���?��)��)�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?G���w��?�B�I .�?�������?�������?_�_��?�A�A�?              �?      �?        .�jL��?IT�n��?ى�؉��?;�;��?�������?UUUUUU�?      �?      �?      �?      �?      �?                      �?      �?              �?                      �?j�V���?Y�����?333333�?�������?              �?�.�袋�?F]t�E�?�������?�������?              �?      �?              �?        �#�;��?w�qGܡ?��<��<�?�a�a�?1P�M��?��k���?��y��y�?�a�a�?      �?              �?      �?              �?      �?              �?                      �?      �?      �?      �?                      �?r�q��?�q�q�?              �?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?              �?      �?      �?              �?      �?              �?      �?        �������?ZZZZZZ�?              �?�������?UUUUUU�?�?�?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?      �?              �?      �?        \�9	ą�?�+c���?	�%����?{	�%���?�q�q�?9��8���?      �?      �?;�;��?�؉�؉�?UUUUUU�?�������?      �?      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?              �?      �?      �?      �?                      �?      �?      �?              �?      �?              �?      �?              �?      �?        �`�`�?�>�>��?�;�;�?�؉�؉�?�������?333333�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?              �?              �?      �?        �k(���?(�����?      �?        333333�?�������?              �?      �?        �������?�������?              �?�������?�������?9��8���?�q�q�?              �?      �?                      �?)M�|�?��,����?     ��?      �?e�M6�d�?N6�d�M�?      �?      �?ffffff�?333333�?              �?9��8���?�q�q�?              �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?^Cy�5�?(������?      �?      �?      �?                      �?              �?�{����?�B!��?�m۶m��?�$I�$I�?      �?        �5��P�?(�����?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?���fy�?�Y�D�a�?߫�^H�?U{���?�ˠT�?ޏ��k��?����v��?�O�%�L�?�RJ)���?[k���Z�?�m۶m��?%I�$I��?�������?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?Y�B��?���7���?�}A_Ч?�/����?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�4��g�?kyc��?qG�wĭ?�;⎸#�?�a�a�?��y��y�?�؉�؉�?��N��N�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?              �?      �?                      �?���k��?7�A�0��?              �?��k���?�@	o4u�?�?�������?              �?�������?�������?              �?      �?        �?�?              �?;�;��?�؉�؉�?      �?                      �?���Q��?)\���(�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?      �?                      �?KԮD�J�?ە�]���?y�5���?�5��P�?      �?        �?�������?              �?;�;��?ى�؉��?              �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?                      �?              �?t�E]t�?��.���?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�?�?              �?      �?      �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�8�hhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�,         n       
             �?z��K���?�           ��@              Q                   �b@>{����?           @y@              $                    �?$�Q�\�?�             u@               	                    �?�P��G7�?H            @]@                                   \@�G��l��?             5@        ������������������������       �                     @                                   a@�q�q�?
             .@       ������������������������       �                     $@        ������������������������       �                     @        
              
             �?��8����?:             X@                                  @_@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @               #       	          ����?���W���?6            �U@                                 �]@     ��?             H@        ������������������������       �                     *@                                  �_@��R[s�?            �A@                                  `X@      �?             0@                                  @`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             &@               "                    �?D�n�3�?             3@                     	          ����?ҳ�wY;�?             1@                                  �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                      	            �?X�<ݚ�?             "@        ������������������������       �                      @               !                    �?և���X�?             @                                  l@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     C@        %       B                   @^@�IєX�?�            �k@       &       =       	          ����?�7���?Q             _@        '       <                   �`@�����?"            �H@       (       ;                    �?     ��?             @@       )       ,                    �?�4�����?             ?@        *       +                   @Z@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        -       8                   �]@"pc�
�?             6@       .       /       	          ����?R���Q�?             4@       ������������������������       �        	             &@        0       1                    ^@�q�q�?             "@        ������������������������       �                     @        2       3                    `@���Q��?             @        ������������������������       �                     �?        4       5                   �Y@      �?             @        ������������������������       �                     �?        6       7                   l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        9       :                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        >       ?                   �c@�}��L�?/            �R@       ������������������������       �        &            �K@        @       A                    �Q@P���Q�?	             4@       ������������������������       �                     3@        ������������������������       �                     �?        C       N                    f@`�E���?F            @X@       D       M                   `@�L��ȕ?B            @W@        E       L                    �?Pa�	�?            �@@       F       G                   �_@���7�?             6@       ������������������������       �                     3@        H       K       	             �?�q�q�?             @       I       J                   pk@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �        )             N@        O       P                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        R       ]                    �?�\����?,            �P@        S       \                    @��H�}�?             9@       T       U                   �\@���N8�?             5@        ������������������������       �                     �?        V       [       	          ����?z�G�z�?             4@       W       X                   �d@�IєX�?             1@       ������������������������       �                     &@        Y       Z                   �_@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ^       _                    c@��]�T��?            �D@        ������������������������       �                     @        `       a                   �c@�����?             C@        ������������������������       �        
             ,@        b       c                    �?      �?             8@        ������������������������       �                     @        d       i                   �^@p�ݯ��?             3@       e       h                   e@�θ�?             *@        f       g       
             �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        j       m                   �p@�q�q�?             @       k       l                    d@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        o       �       	            �?`m��A�?�            �t@       p       �                    �M@����"$�?�             p@       q       �                    �?~~���?�            �m@        r       }                    �?      �?             L@       s       t                     D@�:�^���?            �F@        ������������������������       �                     (@        u       |                    ]@<���D�?            �@@        v       w                   @[@�q�q�?	             (@        ������������������������       �                      @        x       y                   �b@���Q��?             $@        ������������������������       �                     @        z       {                   d@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        ~                          pq@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        �       �                    �?����?�?f            �f@       �       �                   �l@@��'��?[             d@       ������������������������       �        0            �U@        �       �                    �?��
���?+            �R@        ������������������������       �                     @@        �       �                   `d@ �#�Ѵ�?            �E@       ������������������������       �                     =@        �       �       	          ����?؇���X�?	             ,@       �       �                     J@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        �       �                   �`@�KM�]�?             3@       ������������������������       �                     &@        �       �                   @b@      �?              @        ������������������������       �                     @        �       �                   @a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�eP*L��?             6@       �       �                   xt@r�q��?             (@       �       �                    �N@�C��2(�?             &@        �       �                   xs@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?X�<ݚ�?/             R@       �       �                   �^@��X��?$             L@        ������������������������       �                     "@        �       �                   ``@��k=.��?            �G@        ������������������������       �                     1@        �       �                    �N@�z�G��?             >@       �       �                    b@�û��|�?             7@       �       �       	          ����?�	j*D�?	             *@       �       �                    @L@�q�q�?             @        ������������������������       �                      @        �       �                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        �       �                   �Z@      �?             0@       ������������������������       �                     *@        �       �       	          033�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  K�ۚ��?�)|�� �?3|#
L:�?� w�l��?�	j*D�?)ݾ�z��?��)��)�?Z��Y���?��y��y�?1�0��?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?�������?333333�?              �?      �?        ���)kʺ?*kʚ���?      �?      �?              �?PuPu�?X|�W|��?      �?      �?�������?�������?      �?                      �?              �?(������?l(�����?�������?�������?      �?      �?      �?                      �?r�q��?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?      �?                      �?�?�?��Zk���?)��RJ)�?����X�?^N��)x�?      �?      �?��RJ)��?���Zk��?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?/�袋.�?333333�?333333�?              �?UUUUUU�?UUUUUU�?              �?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?                      �?              �?O贁N�?�_,�Œ�?              �?�������?ffffff�?              �?      �?        ����??��W�?X`��?��~���?|���?|���?F]t�E�?�.�袋�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?              �?      �?      �?      �?                      �?>����?���>��?{�G�z�?
ףp=
�?�a�a�?��y��y�?              �?�������?�������?�?�?      �?        �������?UUUUUU�?              �?      �?                      �?              �?jW�v%j�?KԮD�J�?      �?        ^Cy�5�?Q^Cy��?              �?      �?      �?              �?^Cy�5�?Cy�5��?ى�؉��?�؉�؉�?�$I�$I�?۶m۶m�?              �?      �?              �?        UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?        �
ŭP��?���H���?YS֔5e�?6eMYSִ?���c+��?�A�Iݧ?      �?      �?}�'}�'�?l�l��?      �?        |���?|���?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?        �������?�������?              �?      �?              �?        F]t�E�?t�E]t�?      �?                      �?��I��I�?l�l��?�l<��?r���p�?      �?        &�X�%�?O贁N�?      �?        �/����?�}A_Ч?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?        �k(���?(�����?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        t�E]t�?]t�E�?�������?UUUUUU�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�������?              �?      �?        r�q��?�q�q�?n۶m۶�?%I�$I��?              �?g���Q��?br1���?      �?        ffffff�?333333�?8��Moz�?��,d!�?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJP�dhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@/         v                    �?8}�ý�?�           ��@              C       
             �?�q�q�?           0{@               4                    �?h�n��?e            @e@                                  �F@*;L]n�?B             ^@               
                   �[@�z�G��?             >@                                  Pp@�q�q�?             "@       ������������������������       �                     @               	                   q@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                   @D@؇���X�?
             5@                                  �]@���!pc�?             &@        ������������������������       �                     @                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@               !                    �?P�%f��?3            �V@                                  �c@      �?             8@                                 @a@�r����?
             .@        ������������������������       �                     "@                                   �?�q�q�?             @                                  @O@�q�q�?             @                     
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                       	          ����?�<ݚ�?             "@                                 �o@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        "       3                   `c@r٣����?&            �P@       #       $                    �J@Z���c��?$            �O@        ������������������������       �                     5@        %       .       	          @33�?��i#[�?             E@        &       +                    �?���Q��?             4@        '       (       	          ����?X�<ݚ�?             "@        ������������������������       �                     @        )       *                   �b@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ,       -                    �K@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        /       0                    @O@���7�?             6@       ������������������������       �                     0@        1       2                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        5       >                   �b@H%u��?#             I@       6       ;                    @������?            �D@       7       :                    @M@������?             B@        8       9                   8w@�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?        ������������������������       �                     3@        <       =                    `P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       @                   `@X�<ݚ�?             "@        ������������������������       �                     @        A       B                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        D       u       	          ���@pe����?�            �p@       E       X                    @L@�]�{���?�            0p@       F       K                    @H@�}�+r��?�             j@       G       J                    �?0�ޤ��?O            @`@        H       I                   �d@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �        D            �]@        L       Q                   �]@$��$�L�?8            �S@        M       N                   �[@և���X�?	             ,@       ������������������������       �                     @        O       P                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        R       W       	             �?��ɉ�?/            @P@       S       T       	          ����?     ��?.             P@       ������������������������       �        +             N@        U       V                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        Y       d                   �b@`�Q��?              I@       Z       a                   P`@д>��C�?             =@        [       ^                    �?X�<ݚ�?             "@       \       ]                    �M@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        _       `                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        b       c                   �V@P���Q�?
             4@        ������������������������       �                     �?        ������������������������       �        	             3@        e       p                   Pd@�G��l��?             5@       f       g                   �g@����X�?
             ,@        ������������������������       �                     �?        h       k                   ``@�θ�?	             *@        i       j                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       m                    �N@ףp=
�?             $@       ������������������������       �                      @        n       o       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        q       t                    �L@؇���X�?             @        r       s                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        w       z                    Z@�,t�r�?�            �r@        x       y                   �m@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        {       �                    �?��1���?�             r@        |       �       	          ����?�99lMt�?            �C@        }       ~                    �?������?
             1@        ������������������������       �                     "@               �       	          ����?      �?              @       �       �                    f@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �G@���7�?             6@        �       �                   0p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        �       �                   �[@ �_�x�?�            `o@        �       �                    �?�q�q�?             5@       �       �                   `_@      �?             (@        ������������������������       �                     @        �       �       	          `ff�?�q�q�?             "@       �       �                     E@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �Z@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?���.�6�?�            �l@       �       �       	          ����?�==Q�P�?u            �g@       �       �                   �_@���N8�?=            @Z@       ������������������������       �        &             N@        �       �       	          ����?�����H�?            �F@       �       �                   pb@�FVQ&�?            �@@       ������������������������       �                     <@        �       �       	          ����?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    b@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        �       �                    �R@`��>�ϗ?8            @U@       ������������������������       �        6            �T@        �       �                   �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �`@R���Q�?             D@        �       �                   q@b�2�tk�?             2@       �       �                   �[@     ��?
             0@        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                   �]@X�<ݚ�?             "@        �       �       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   pf@�C��2(�?             6@       �       �                   �d@���N8�?             5@       ������������������������       �        	             1@        �       �                     K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  a[ӿc�?PR Np�?UUUUUU�?UUUUUU�?�������?�?�������?""""""�?ffffff�?333333�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?F]t�E�?t�E]t�?      �?              �?      �?              �?      �?              �?        �`�`�?�O��O��?      �?      �?�������?�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �q�q�?9��8���?�������?333333�?              �?      �?                      �?|���?>���>�?��i��i�?Y�eY�e�?              �?�<��<��?�a�a�?333333�?�������?�q�q�?r�q��?              �?�������?�������?              �?      �?        F]t�E�?t�E]t�?              �?      �?        F]t�E�?�.�袋�?              �?UUUUUU�?�������?              �?      �?              �?        ���Q��?)\���(�?������?p>�cp�?�q�q�?�q�q�?�?�?              �?      �?                      �?�������?�������?              �?      �?        �q�q�?r�q��?              �?�������?�������?              �?      �?        ��8��?r�8�?�����?��q/�?�5��P�?(�����?/�B/�B�?z�z��?      �?      �?              �?      �?              �?        ��]-n��?�3���?�$I�$I�?۶m۶m�?      �?        �$I�$I�?۶m۶m�?              �?      �?        ?�?��? �����?     ��?      �?      �?              �?      �?              �?      �?                      �?��(\���?{�G�z�?a���{�?|a���?r�q��?�q�q�?�������?�������?              �?      �?              �?      �?      �?                      �?ffffff�?�������?              �?      �?        ��y��y�?1�0��?�$I�$I�?�m۶m��?      �?        �؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?                      �?�C����?/� }J�?�q�q�?�q�q�?      �?                      �?x��ǿ?�p���?�o��o��?5H�4H��?xxxxxx�?�?      �?              �?      �?�������?�������?              �?      �?              �?        F]t�E�?�.�袋�?UUUUUU�?UUUUUU�?      �?                      �?              �?����0p�?g��1�?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?�q�q�?�q�q�?              �?      �?        Y�B��?���7���?�a�+�?��%N��?�a�a�?��y��y�?              �?�q�q�?�q�q�?|���?>����?              �?�������?333333�?              �?      �?              �?      �?              �?      �?        �?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?9��8���?�8��8��?      �?      �?              �?�������?�������?r�q��?�q�q�?�������?�������?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?              �?      �?        F]t�E�?]t�E�?�a�a�?��y��y�?              �?      �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�g?BhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKۅ�h��B�6         |                    �?2��ή�?�           ��@              =                    @L@"` Y��?           �z@              "                    �?h�eX��?�            �q@                      
             �?�q���?=             X@                                  `p@$�q-�?            �C@       ������������������������       �                     <@                      	          ����?���!pc�?             &@        ������������������������       �                     @        	       
                   ``@���Q��?             @        ������������������������       �                     �?                                  Pc@      �?             @        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  `]@P̏����?"            �L@                                  `m@����X�?	             ,@                                 �`@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@                                   �?      �?             @                                 �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?�ʈD��?            �E@                                 �d@P���Q�?             D@       ������������������������       �                     >@                                   e@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @                !                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        #       (                   `R@�_�����?x             g@        $       '                   �^@�q�q�?             "@        %       &                   �K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        )       <       
             �?p}"����?r            �e@        *       +                    �?�G�z�?             D@        ������������������������       �                     &@        ,       ;                    �?П[;U��?             =@       -       2                    �G@r�q��?             8@        .       /                   �m@���!pc�?             &@       ������������������������       �                     @        0       1                   �r@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        3       8                    �?�θ�?	             *@        4       7                   �c@�q�q�?             @       5       6                   @q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        9       :                    \@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �        Y            �`@        >       _       
             �?��Q����?W            @b@       ?       D                   `\@*�s���?2             U@        @       C                   `Q@�}�+r��?             C@        A       B                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     A@        E       J                   `@�I� �?             G@        F       I                    l@�q�q�?             (@       G       H       	             �?���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        K       P                   `k@H�V�e��?             A@       L       M       	          ���@P���Q�?             4@       ������������������������       �        	             *@        N       O                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        Q       X                    �M@և���X�?             ,@        R       S                   c@�q�q�?             @        ������������������������       �                     @        T       U                   d@�q�q�?             @        ������������������������       �                     �?        V       W                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                    �?      �?              @        ������������������������       �                     @        [       \                    �?      �?             @        ������������������������       �                     �?        ]       ^                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        `       {       	          ���@�4�����?%             O@       a       z                   @e@�c�Α�?"             M@       b       g                   �V@�\�u��?            �I@        c       d       	          ���ɿ���Q��?             $@        ������������������������       �                      @        e       f                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        h       u                    s@���?            �D@       i       t                    �N@     ��?             @@        j       q       	          ����?X�Cc�?	             ,@       k       l                    d@z�G�z�?             $@        ������������������������       �                     @        m       n                    �L@�q�q�?             @        ������������������������       �                     �?        o       p                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        r       s                   p`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             2@        v       y                   �u@X�<ݚ�?             "@       w       x                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        }       �       
             �?�䞠�l�?�            @s@       ~       �                    @�L���?�            0p@              �                    �?     ��?�             p@       �       �                   @b@������?�             j@       �       �       	          033�?�O���h�?|            �f@        �       �                    �?��p\�?            �D@       �       �                    f@      �?             8@       �       �       	          ����?���}<S�?             7@       ������������������������       �                     0@        �       �       	          hff�?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             1@        �       �                   @X@@P���x�?b            �a@        �       �                   �`@�C��2(�?             &@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �_@ g�yB�?Z             `@       �       �                   `_@�(\����?8             T@       �       �                   �r@`׀�:M�?3            �R@       ������������������������       �        *             N@        �       �                    �Q@@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        �       �       	          ����?r�q��?             @        ������������������������       �                      @        �       �                   �j@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        "            �H@        �       �                    �?�+$�jP�?             ;@       �       �                   pn@�q�q�?	             .@        �       �                   �h@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     (@        �       �                    @G@8��8���?!             H@        ������������������������       �                      @        �       �                    �?�q��/��?             G@        �       �       	             �?z�G�z�?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@������?            �D@       �       �                   �\@ >�֕�?            �A@        �       �       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @^@      �?             @@        �       �                   Xr@@4և���?
             ,@       ������������������������       �                     (@        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             2@        �       �                     M@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �I@~���L0�?            �H@        �       �                   pq@X�Cc�?	             ,@       �       �                   �Z@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                   �e@b�h�d.�?            �A@       �       �                   �`@��hJ,�?             A@       �       �                    �?�C��2(�?             6@       �       �                   �^@�IєX�?             1@        �       �                    �?؇���X�?             @        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    _@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �`@      �?
             (@        ������������������������       �                     �?        �       �                   �a@"pc�
�?	             &@        ������������������������       �                     @        �       �       	          ����?����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  7�@c��?d�_yΨ�?�V�H�?��RO�o�?�A�A�?�������?�������?�������?;�;��?�؉�؉�?              �?t�E]t�?F]t�E�?              �?333333�?�������?              �?      �?      �?      �?              �?      �?              �?      �?        ?���#�?��Gp�?�$I�$I�?�m۶m��?�������?�������?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        A_���?�}A_з?ffffff�?�������?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        Y�B��?�7��Mo�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?ĦҐs��?��jyc�?�������?�������?      �?        �{a���?��=���?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?      �?              �?      �?              �?      �?        �؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �������?�������?      �?                      �?      �?              �?        ϝ;w���?1bĈ�?z��y���?b�a��?(�����?�5��P�?      �?      �?      �?                      �?              �?Nozӛ��?Y�B���?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?              �?      �?                      �?ZZZZZZ�?iiiiii�?�������?ffffff�?              �?�$I�$I�?۶m۶m�?              �?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?���Zk��?��RJ)��?5�rO#,�?�{a���?�������?�?�������?333333�?      �?              �?      �?      �?                      �?28��1�?8��18�?      �?      �?%I�$I��?�m۶m��?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?              �?      �?              �?        �q�q�?r�q��?UUUUUU�?�������?              �?      �?              �?              �?                      �?5�wL�?�	qV~B�?L�Ϻ��?}���g�?      �?     ��?;�;��?��N��N�?������?�0&q��?��+Q��?�]�ڕ��?      �?      �?d!Y�B�?ӛ���7�?              �?�$I�$I�?�m۶m��?      �?                      �?      �?                      �?_�_�?uPuP�?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?����?�����?�������?333333�?к����?��L��?              �?�$I�$I�?n۶m۶�?              �?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?B{	�%��?/�����?UUUUUU�?UUUUUU�?�������?UUUUUU�?              �?      �?                      �?              �?�������?UUUUUU�?      �?        ��Mozӻ?�B����?�������?�������?              �?      �?      �?      �?                      �?������?�|����?�A�A�?��+��+�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        ������?����>4�?%I�$I��?�m۶m��?�������?�������?              �?      �?                      �?_�_��?;��:���?�������?KKKKKK�?F]t�E�?]t�E�?�?�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�������?              �?      �?              �?      �?      �?        F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ1�.hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKǅ�h��B�1         v                    �?�������?�           ��@              Q                    �?��Q����?           Py@                                  �?x9G����?�            �s@                      	          `ff�?�̐d��?I            @Z@                                  �?p�|�i�?6             S@                                  �b@      �?             (@        ������������������������       �                     @                                  �b@      �?              @       	       
       
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        .             P@                      
             �?J�8���?             =@                                  b@�G��l��?             5@                                 p@r�q��?	             (@       ������������������������       �                      @                                   �?      �?             @        ������������������������       �                     �?                      	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                      
             �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               <       
             �?8�Z$(�?�             j@                                  `\@�A����?6            �T@        ������������������������       �        	             ,@                                  @^@.Lj���?-             Q@        ������������������������       �                     @                -                    @J@�	j*D�?*            @P@       !       ,                   �`@     ��?             @@       "       +                   `r@�����?             3@       #       &                    �?������?             1@        $       %                   8p@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        '       (                    �?�8��8��?             (@        ������������������������       �                     @        )       *                   @g@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        .       9       	          pff�?4���C�?            �@@       /       0                   �_@�E��ӭ�?
             2@        ������������������������       �                     "@        1       8                   Pp@X�<ݚ�?             "@       2       7                   @k@և���X�?             @       3       6                   Pi@      �?             @       4       5                   a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        :       ;                   �d@��S�ۿ?	             .@       ������������������������       �                     ,@        ������������������������       �                     �?        =       H       	          ����?�����H�?Q            �_@       >       G                   �t@`�q�0ܴ?=            �W@       ?       F                   0m@��<b�ƥ?<             W@       @       E                   �l@`2U0*��?!             I@       A       B                    b@@�E�x�?             �H@       ������������������������       �                    �B@        C       D                   �b@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     E@        ������������������������       �                      @        I       P                    �?     ��?             @@       J       K                   @a@��}*_��?             ;@        ������������������������       �                     @        L       M                    @K@�G��l��?             5@        ������������������������       �                     @        N       O       	          ����?�q�q�?             .@        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @        R       [                    �?�I� �?4             W@        S       Z                   �c@"pc�
�?             &@       T       Y                    �?�q�q�?             @       U       X                    �?�q�q�?             @       V       W                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        \       a                   �`@������?.            @T@        ]       ^                    @��<b�ƥ?             G@       ������������������������       �                     C@        _       `                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        b       u       	          ���	@և���X�?            �A@       c       d                    �E@      �?             @@        ������������������������       �                     @        e       n                    �M@������?             ;@       f       i                    �?��s����?             5@        g       h       
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        j       k                    �?�IєX�?             1@       ������������������������       �        	             ,@        l       m                   @^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        o       p                   �`@      �?             @        ������������������������       �                      @        q       r                   �V@      �?             @        ������������������������       �                      @        s       t                    �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        w       �                    �?��E�B��?�            �t@       x       �                    �?̘#ZJ�?�            �p@        y       z                    m@4�2%ޑ�?            �A@        ������������������������       �                     (@        {       |       	          ����?�LQ�1	�?             7@        ������������������������       �                     @        }       �                    @I@�t����?             1@        ~                          �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@��S�ۿ?	             .@        �       �       	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                   �d@���.�6�?�            �l@       �       �                    `R@�yr�?c�?�            �l@       �       �                    �? '��h�?�            @k@       �       �                   �[@���C�:�?_            `b@        �       �                   ph@X�<ݚ�?             "@        ������������������������       �                      @        �       �       	             �?և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   0q@�nkK�?X            @a@       �       �                    q@0G���ջ?C             Z@       �       �       
             �?X�?٥�?B            �Y@       �       �                    \@F|/ߨ�?4            @T@        �       �                   p@@-�_ .�?            �B@       ������������������������       �                     @@        �       �                    Z@���Q��?             @        ������������������������       �                      @        �       �                   �_@�q�q�?             @       �       �                   pp@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     F@        �       �                    c@��2(&�?             6@       �       �                    �I@P���Q�?             4@        �       �                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             0@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     A@        ������������������������       �        ,            �Q@        �       �       
             �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @     ��?%             P@       �       �                   �`@�&�5y�?$             O@       �       �       
             �?t��ճC�?             F@       �       �                   P`@�Ń��̧?             E@        �       �                     N@��S�ۿ?
             .@        �       �                    �L@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@        ������������������������       �                      @        �       �                   ``@�<ݚ�?             2@        �       �                   �[@      �?             @        ������������������������       �                      @        �       �       
             �?      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�8��8��?             (@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  -@��"�?�߱����?;��WaN�?��FP=c�?b�c�)5�?<o8����?��	��	�? �����?�k(����?^Cy�5�?      �?      �?      �?              �?      �?�������?UUUUUU�?              �?      �?                      �?      �?        �rO#,��?|a���?1�0��?��y��y�?�������?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?      �?                      �?      �?        O��N���?b'vb'v�?�18���?�cp>�?              �?�������?------�?      �?        ;�;��?vb'vb'�?      �?      �?^Cy�5�?Q^Cy��?�?xxxxxx�?333333�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?'�l��&�?m��&�l�?�q�q�?r�q��?      �?        �q�q�?r�q��?�$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?�?�������?              �?      �?        �q�q�?�q�q�?��F}g��?W�+�ɥ?��7��M�?d!Y�B�?���Q��?{�G�z�?և���X�?9/���?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?      �?_B{	�%�?B{	�%��?      �?        1�0��?��y��y�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        Nozӛ��?Y�B���?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?              �?        {	�%���?B{	�%��?d!Y�B�?��7��M�?              �?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?B{	�%��?{	�%���?z��y���?�a�a�?      �?      �?              �?      �?        �?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?              �?      �?              �?      �?      �?              �?      �?                      �?AL� &W�?�l�w6��?�q�8�?>���8�?�A�A�?�������?              �?d!Y�B�?Nozӛ��?      �?        �?<<<<<<�?      �?      �?      �?                      �?�?�������?      �?      �?      �?                      �?              �?Y�B��?���7���?˂��"M�?���-�?�w� z|�?���]8��?[��5;j�?uo@����?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?d!Y�B�?�Mozӛ�?�؉�؉�?vb'vb'�?C��ڨ?�">�Tr�?�����H�?�Hx�5�?к����?S�n0E�?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?t�E]t�?��.���?�������?ffffff�?      �?      �?      �?                      �?              �?      �?              �?                      �?              �?F]t�E�?]t�E]�?      �?                      �?      �?              �?     ��?�1�c��?:�s�9�?t�E]t�?�E]t��?�a�a�?��<��<�?�?�������?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?      �?        9��8���?�q�q�?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �t�bub��     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJg�)hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKم�h��B@6         ~                    �?$~��,��?�           ��@              -                    �J@������?�            Py@                                   �?�npº��?[            �b@                                   �?      �?*             T@                                 Hq@�t����?!             Q@              	       
             �?��f/w�?            �N@                                  �p@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        
                           �I@@��8��?             H@       ������������������������       �                     E@                                   m@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   @H@r�q��?	             (@        ������������������������       �                     @                                  �]@�q�q�?             @                                  ]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               ,                   pf@D��\��?1            �Q@                                 �Z@������?0            �Q@        ������������������������       �                      @                                  �[@ДX��?/             Q@                                  �`@����X�?             @       ������������������������       �                     @                      	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                +                   �p@85�}C�?*            �N@       !       &                    �?6YE�t�?            �@@        "       #                   �\@և���X�?             @        ������������������������       �                      @        $       %                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        '       (       	             @$�q-�?             :@       ������������������������       �                     6@        )       *                   �o@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     <@        ������������������������       �                     �?        .       U                    �?Po��ب�?�            �o@        /       T                   �c@���%&�?0            �S@       0       I       	          ����?�Jhu4��?+            @R@       1       D                   Pc@\X��t�?             G@       2       7                   @E@<ݚ)�?             B@        3       4       	             �?      �?              @       ������������������������       �                     @        5       6                   �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        8       C       
             �?�>4և��?             <@       9       @                    �?     ��?	             0@       :       ?                   �_@�θ�?             *@       ;       <                    �?      �?             @        ������������������������       �                     �?        =       >                   �q@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        A       B       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        E       F                   �`@ףp=
�?             $@        ������������������������       �                     @        G       H                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        J       S       	             �?PN��T'�?             ;@        K       R                    �?����X�?             ,@       L       Q                    �P@�θ�?             *@       M       N                    c@r�q��?             (@       ������������������������       �                     "@        O       P                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     @        V       y                    c@�#-���?s            �e@       W       x       	          ��� @@4և���?m             e@       X       m                   (r@\#r��?S            �^@       Y       b                   `_@0G���ջ?F             Z@       Z       a                    �?�(\����?3             T@       [       `                   �[@ �q�q�?             H@       \       _                    �L@�>����?             ;@        ]       ^                   pm@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     6@        ������������������������       �                     5@        ������������������������       �                     @@        c       j                   @U@r�q��?             8@        d       e       
             �?և���X�?             @        ������������������������       �                     @        f       i                   �`@      �?             @       g       h                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        k       l                   @]@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �                     0@        n       s       	          ����?�q�q�?             2@        o       p       	          ����?r�q��?             @        ������������������������       �                     @        q       r                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        t       u                    c@�8��8��?	             (@       ������������������������       �                     $@        v       w                    `P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     G@        z       }                    q@և���X�?             @       {       |                   �d@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               �       
             �?�����?�            �t@        �       �                    �?"` Y��?W            �a@        �       �                   xu@�θ�?             :@       �       �                   �b@r�q��?             8@       �       �                   �Q@�LQ�1	�?             7@        ������������������������       �                     �?        �       �                   �Z@�C��2(�?             6@        ������������������������       �                     �?        �       �                   �e@���N8�?             5@       ������������������������       �                     1@        �       �                    �I@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   a@�c�Α�?D             ]@       �       �       
             �?85�}C�?$            �N@        �       �                    �?�q�q�?             @        �       �                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     F@�1�`jg�?             �K@        �       �                   @_@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?`2U0*��?             I@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @L@����?�?            �F@        �       �                   `_@�C��2(�?             &@        �       �                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     A@        �       �                   b@D7�J��?             �K@        �       �                   �a@     ��?	             0@       �       �                   �a@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �m@�e����?            �C@       �       �                   m@R�}e�.�?             :@       �       �                   �^@�q�q�?             5@        ������������������������       �                     @        �       �                    @N@��S���?
             .@       �       �                    _@      �?              @        ������������������������       �                     �?        �       �                     F@؇���X�?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          pff�?�	j*D�?	             *@       ������������������������       �                     "@        ������������������������       �                     @        �       �                    �? ��@��?~            `g@       �       �       	          ���@8�Z� �?n            `d@       �       �                    @L@�fp�IЮ?l             d@       �       �                   �_@ �|ك�?R            �^@        �       �                   �^@�8��8��?             (@       ������������������������       �        
             &@        ������������������������       �                     �?        ������������������������       �        G            �[@        �       �                    �M@�KM�]�?             C@        �       �                   �r@�<ݚ�?             2@       �       �                    d@�r����?
             .@        ������������������������       �                     @        �       �                    a@      �?              @        ������������������������       �                     �?        �       �                    c@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                      @        �       �                   �U@      �?             8@        �       �       	          ����?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��C�l��??+^�ɑ�?{	�%���?B{	�%��?˸e�2n�?�#͑�H�?      �?      �?�������?�������?XG��).�?��!XG�?;�;��?�؉�؉�?              �?      �?        UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?              �?      �?                      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?�@�6�?�o�z2~�?PuPu�?,��+���?      �?        ZZZZZZ�?�������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        ������?�}�K�`�?e�M6�d�?'�l��&�?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?;�;��?�؉�؉�?              �?      �?      �?              �?      �?                      �?      �?        ��j�Z��?�J�R�T�?�0���M�?�g *��?ҤI�&M�?�-[�l��?!Y�B�?��Moz��?��8��8�?�8��8��?      �?      �?              �?      �?      �?              �?      �?        �$I�$I�?�m۶m��?      �?      �?ى�؉��?�؉�؉�?      �?      �?      �?        �������?333333�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?h/�����?&���^B�?�$I�$I�?�m۶m��?�؉�؉�?ى�؉��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?              �?_�_�?�A�A�?�$I�$I�?n۶m۶�?XG��).�?��:��?�؉�؉�?vb'vb'�?�������?333333�?UUUUUU�?�������?h/�����?�Kh/��?�������?333333�?      �?                      �?              �?              �?              �?UUUUUU�?�������?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?              �?      �?              �?        �?�?      �?                      �?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?        ���T��?u�^V	�?��RO�o�?�V�H�?ى�؉��?�؉�؉�?�������?UUUUUU�?��Moz��?Y�B��?              �?]t�E�?F]t�E�?              �?��y��y�?�a�a�?      �?              �?      �?      �?                      �?              �?              �?�{a���?5�rO#,�?������?�}�K�`�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?�־a�?A��)A�?�������?�������?              �?      �?        {�G�z�?���Q��?�������?�������?              �?      �?      �?              �?      �?        l�l��?��I��I�?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?              �?k߰�k�?J��yJ�?      �?      �?      �?      �?              �?      �?              �?        �A�A�?�-��-��?�;�;�?'vb'vb�?UUUUUU�?UUUUUU�?              �?�������?�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?�m۶m��?�$I�$I�?              �?      �?                      �?vb'vb'�?;�;��?      �?                      �?��:����?�)��˱?���A2��?�Ŗ����?̀O��?��6͟?�_��e��?�h
���?UUUUUU�?UUUUUU�?      �?                      �?      �?        �k(���?(�����?9��8���?�q�q�?�������?�?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�]_AhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         R                    @K@znt��s�?�           ��@               )       	          ����?��U�?�            �v@              
                   �Q@��a̒�?�             m@                      
             �?�n`���?             ?@       ������������������������       �                     2@               	       	          ����?��
ц��?             *@                                  �?�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               "                    �?t(d��?~            @i@              !                   �`@��`ۻ��?s            �g@                     
             �?��27
��?U            `a@                                  q@     ��?             @@                     	          ����?l��
I��?             ;@                                   F@���!pc�?             &@        ������������������������       �                     �?                                  �`@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     @                                   `\@�r�MȢ?D            �Z@                                   �?@4և���?             <@                                  c@�q�q�?             @        ������������������������       �                     @                                  �[@�q�q�?             @                                 �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �        1            �S@        ������������������������       �                    �H@        #       (       	          ����?����X�?             ,@       $       %       
             �?r�q��?
             (@       ������������������������       �                      @        &       '                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        *       A                    �?DpJ��?O            ``@        +       8       	          033�?r�q��?             H@        ,       3                   @_@���!pc�?             6@        -       0                   `]@�eP*L��?             &@       .       /       
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        1       2                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        4       7                    �?�C��2(�?             &@        5       6       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        9       :                   �`@�n_Y�K�?             :@        ������������������������       �                     &@        ;       <                   0d@�q�q�?	             .@        ������������������������       �                     @        =       @                   b@r�q��?             (@        >       ?                   pf@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        B       K                   �c@��`qM|�?2            �T@       C       F                   �Z@ ���J��?.            �S@        D       E                   �Y@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        G       J                    \@�}��L�?+            �R@        H       I                   �[@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �        #             O@        L       M       
             �?���Q��?             @        ������������������������       �                     �?        N       O       	          ����?      �?             @        ������������������������       �                      @        P       Q                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       �                    �?�a��+*�?�             w@       T       �       
             �?�c����?�             k@       U       ~                    �?��CC`)�?|            �f@       V       k                   ``@>4և�z�?N             \@        W       X       	          ����?����X�?             E@        ������������������������       �        	             ,@        Y       f                    �?և���X�?             <@       Z       _       	          ����?�d�����?             3@        [       \                    �?z�G�z�?             @        ������������������������       �                     @        ]       ^                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        `       a                    �?@4և���?
             ,@       ������������������������       �                     $@        b       e       	          `ff�?      �?             @        c       d                    ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        g       h                    @L@�<ݚ�?             "@        ������������������������       �                     �?        i       j       	             @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        l       }                    @O@@4և���?1            �Q@       m       v       	          ����?      �?             D@        n       u                   xs@      �?              @       o       t                   �[@����X�?             @       p       s                    b@      �?             @       q       r                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        w       x                    c@      �?             @@       ������������������������       �                     :@        y       |       	          033�?�q�q�?             @       z       {                   xu@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@               �                   �Q@�nkK�?.            @Q@        �       �       	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?����e��?,            �P@        �       �                   �r@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �        #            �J@        �       �                    �?b�2�tk�?             B@        �       �       	          ����?�8��8��?             (@        �       �                   P`@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @E@r�q��?             8@        �       �                    �?      �?              @       ������������������������       �                     @        �       �                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?
             0@        ������������������������       �                     @        �       �                   b@���|���?             &@       ������������������������       �                     @        �       �                    ]@z�G�z�?             @        ������������������������       �                      @        �       �                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �`@��.k���?V             c@        �       �                    �L@���!pc�?             �K@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                    @P@��k=.��?            �G@       �       �       
             �?(;L]n�?             >@       ������������������������       �                     =@        ������������������������       �                     �?        �       �                    @��.k���?             1@       �       �                    �?X�Cc�?	             ,@        ������������������������       �                     @        �       �                    �?"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        �       �       
             �?4=�%�?6            �X@       �       �                   hq@�E��
��?             J@       �       �                   �m@��%��?            �B@       �       �                    �?
j*D>�?             :@        ������������������������       �                     @        �       �                    d@
;&����?             7@       �       �                    �N@p�ݯ��?             3@       �       �                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?؇���X�?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �b@"pc�
�?             &@       �       �                     P@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   Pr@��S�ۿ?             .@       ������������������������       �                     $@        �       �                    �K@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          `ff�?��<b���?             G@       �       �                   �s@,���i�?            �D@       �       �                   �i@      �?             @@        �       �                    d@�����H�?             "@       ������������������������       �                     @        �       �                     M@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                   u@X�<ݚ�?             "@       �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  ����?��}t��?�������?˨�ʨ��?{�a"�?��x�w�?�c�1��?�9�s��?              �?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?      �?                      �?              �?m�2|#
�?�tj䮿?��
br�?R�٨�l�?�j����?p�l�:��?      �?      �?Lh/����?h/�����?t�E]t�?F]t�E�?      �?        �������?�������?              �?      �?              �?                      �?z����f�?�+J�#�?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?              �?              �?        �$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?        J�eDP�?m��.���?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?t�E]t�?]t�E�?�������?UUUUUU�?              �?      �?        �������?�������?              �?      �?        ]t�E�?F]t�E�?      �?      �?              �?      �?              �?        ى�؉��?;�;��?              �?UUUUUU�?UUUUUU�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        ��k���?�@	o4u�?�A�A�?��-��-�?UUUUUU�?UUUUUU�?              �?      �?        O贁N�?�_,�Œ�?;�;��?�؉�؉�?              �?      �?                      �?�������?333333�?      �?              �?      �?              �?      �?      �?      �?                      �?]%�j�U�?Rm�J��?�8P(�?����u��?4O��I�?�J�v�?۶m۶m�?I�$I�$�?�$I�$I�?�m۶m��?              �?۶m۶m�?�$I�$I�?y�5���?Cy�5��?�������?�������?      �?              �?      �?      �?                      �?�$I�$I�?n۶m۶�?              �?      �?      �?      �?      �?              �?      �?                      �?9��8���?�q�q�?              �?      �?      �?      �?                      �?�$I�$I�?n۶m۶�?      �?      �?      �?      �?�$I�$I�?�m۶m��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?d!Y�B�?�Mozӛ�?UUUUUU�?UUUUUU�?              �?      �?        |���?�>����?;�;��?�؉�؉�?              �?      �?                      �?9��8���?�8��8��?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?              �?      �?              �?      �?      �?        ]t�E]�?F]t�E�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �?�������?t�E]t�?F]t�E�?      �?      �?      �?                      �?br1���?g���Q��?�?�������?              �?      �?        �?�������?�m۶m��?%I�$I��?      �?        F]t�E�?/�袋.�?      �?                      �?      �?        ������?�>4և��?��؉���?;�;��?���L�?}���g�?;�;��?b'vb'v�?              �?�Mozӛ�?Y�B��?Cy�5��?^Cy�5�?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?              �?        /�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �?�������?              �?�������?�������?              �?      �?        ��,d!�?��Moz��?�����?8��18�?      �?      �?�q�q�?�q�q�?      �?              �?      �?      �?                      �?      �?        r�q��?�q�q�?�������?�������?              �?      �?      �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJL�OhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         �       
             �?���:���?�           ��@              o       	          ����?ęI0�?           pz@                                 �c@��CU�q�?�            �q@                                   �?�ȉo(��?9            �V@                                  �c@���}<S�?             G@                                 �d@ �#�Ѵ�?            �E@                                  �?��Y��]�?            �D@                                   �?      �?             0@       	       
                   �^@�8��8��?             (@        ������������������������       �                     @                                    O@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@                      	          @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �F@               D                    �?��˹f�?�             h@               '                    �?>����?<            �X@               $                   �r@<ݚ)�?             B@                                 �]@؇���X�?             <@        ������������������������       �                     &@                                   �?������?             1@        ������������������������       �                      @               #                   pd@�r����?             .@                                   �J@      �?              @        ������������������������       �                     @        !       "                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        %       &                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        (       ?                    �?b����?&            �O@       )       *                   `X@����X�?              L@        ������������������������       �                     @        +       8                   hq@�c�����?            �J@       ,       -                    m@���V��?            �F@        ������������������������       �                     3@        .       3                    �?R�}e�.�?             :@       /       2                   �m@8�Z$���?             *@        0       1                   �e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        4       7                     J@�n_Y�K�?             *@        5       6       	          pff�?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        9       <                     @      �?              @       :       ;                   @`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        =       >                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        @       C                    `@؇���X�?             @        A       B                     Q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        E       \                    �?�9�a��?E            �W@       F       W                    �?�θV�?6            @Q@       G       T                    �O@�q��/��?(            �H@       H       I                   `_@�q��/��?%             G@       ������������������������       �                     7@        J       K                   Pf@��<b���?             7@        ������������������������       �                      @        L       O                   �\@؇���X�?             5@        M       N                   @a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        P       S                    �?      �?             0@        Q       R       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        U       V                    o@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        X       [                    Z@P���Q�?             4@        Y       Z                   (q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ]       j       	          ����?���Q��?             9@       ^       _                   j@��.k���?             1@        ������������������������       �                     @        `       e                   �l@�n_Y�K�?	             *@        a       b                   �\@؇���X�?             @        ������������������������       �                     @        c       d       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        f       i                   �a@�q�q�?             @       g       h                    @M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        k       l                    @      �?              @        ������������������������       �                     @        m       n                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        p       s                     E@���۟�?V            `a@        q       r                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        t       �       	          `ff@�����?T            �`@       u       �                     R@ ,V�ނ�?O            �_@       v                          `b@ ��+,��?N            @_@       w       ~                    �?�H�I���?D            @\@       x       y                   8p@�eGk�T�?9            �W@       ������������������������       �        '             O@        z       {       	          033@Pa�	�?            �@@       ������������������������       �                     4@        |       }                    �J@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     2@        �       �                   �q@      �?
             (@       �       �                   �i@      �?             @        ������������������������       �                      @        �       �                   `d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    P@4�Q�]�?�            ps@        �       �                    �?h+�v:�?             A@       �       �                    �?      �?             8@       �       �                    �?     ��?             0@        �       �                   �_@      �?             @        �       �                    �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �       	          @33�?      �?              @        �       �                   �a@      �?             @       �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��e��?�            Pq@        �       �                    �?p���?@             Y@        �       �                    b@؇���X�?	             ,@       ������������������������       �                     $@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        7            �U@        �       �                    �?Z��@�}�?t             f@        �       �                   �a@��7��?,            �N@        �       �                    �L@؇���X�?             <@       ������������������������       �                     5@        �       �                    �?և���X�?             @       �       �       	          ����?z�G�z�?             @        �       �                     O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   `\@4���C�?            �@@        �       �                    �E@�����H�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?r�q��?             8@        �       �                   �i@r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?      �?	             (@        �       �                    o@      �?             @       �       �                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @L@ 	��p�?H             ]@       �       �       	          ����?@�E�x�?;            �X@       ������������������������       �        6             V@        �       �                   �_@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�q�q�?             2@       �       �                   �m@z�G�z�?             $@        �       �                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �a@      �?              @        ������������������������       �                     @        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @`@      �?              @        ������������������������       �                      @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  !��Q��?p��1W-�?�k���?e����?l$Zas�?���RO��?h�h��?�~��?d!Y�B�?ӛ���7�?�}A_Ч?�/����?������?8��18�?      �?      �?UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?)!�~��?ko��@��?z;Cb���?�y;Cb�?�8��8��?��8��8�?�$I�$I�?۶m۶m�?              �?�?xxxxxx�?      �?        �?�������?      �?      �?              �?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?5M�4M��?�eY�eY�?�m۶m��?�$I�$I�?              �?�V�9�&�?:�&oe�?[�[��?�>�>��?      �?        'vb'vb�?�;�;�?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        ;�;��?ى�؉��?�$I�$I�?�m۶m��?              �?      �?              �?              �?      �?UUUUUU�?�������?              �?      �?              �?      �?      �?                      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?]AL� &�?��l�w6�?�Q�g���?̵s���?և���X�?/����?��Mozӻ?�B����?              �?��Moz��?��,d!�?      �?        �$I�$I�?۶m۶m�?�������?333333�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?ffffff�?      �?      �?      �?                      �?              �?�������?333333�?�?�������?              �?;�;��?ى�؉��?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?              �?      �?              �?�������?333333�?      �?                      �?����j�?��a����?�������?�������?              �?      �?        ���@��?g��1��?EQEQ�?�뺮��?����Mb�?`��"���?x�!���?x�!���?�X�0Ҏ�?��=�ĩ�?              �?|���?|���?              �?;�;��?�؉�؉�?      �?                      �?              �?      �?      �?      �?      �?              �?      �?      �?      �?                      �?              �?      �?              �?      �?              �?      �?        ��oH�q�?�4@ޞ9�?xxxxxx�?�������?      �?      �?      �?      �?      �?      �?      �?      �?              �?      �?              �?                      �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?ffffff�?333333�?      �?                      �?�y�0�?�s7���?\���(\�?{�G�z�?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        �,1>e�?ƧL;k�?&C��6��?�y��!�?۶m۶m�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?              �?      �?        '�l��&�?m��&�l�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?�������?UUUUUU�?              �?      �?              �?      �?      �?      �?      �?      �?              �?      �?                      �?              �?������?�{a���?և���X�?9/���?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��lhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKׅ�h��B�5         �                    �?<���m�?�           ��@              k       	          ����?R;;�p`�?           `z@                                 �c@�@���0�?�            �u@                                  �^@���N8�?             E@                                   �?p�ݯ��?             3@                                  �I@r�q��?	             (@                                   �G@      �?             @        ������������������������       �                     �?        	       
                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                   �?����X�?             @                                  �?r�q��?             @        ������������������������       �                     �?                                   @K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                      
             �?�LQ�1	�?             7@                     	            �?�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?                                  `a@���Q��?             @                                 @b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @               D       
             �?���
.��?�            0s@               %                    �F@���%&�?,            �S@               $                   q@�����?             3@               #                   �[@@4և���?	             ,@        !       "                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        &       C                    �?��0u���?              N@       '       :                   0a@�q�q�?            �I@       (       7                   0e@և���X�?            �A@       )       .                   @^@|��?���?             ;@        *       +                    �K@���|���?             &@        ������������������������       �                     @        ,       -       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        /       2                    �?     ��?	             0@       0       1                     M@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        3       4                    �?      �?              @        ������������������������       �                     @        5       6       	          hff�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        8       9                    @H@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ;       <       	          ����?      �?	             0@        ������������������������       �                     @        =       B                    �?z�G�z�?             $@       >       ?                    �N@�����H�?             "@       ������������������������       �                     @        @       A       	          pff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        E       b                   �s@�1Y�I��?�            �l@       F       Y                    �?�V���?�            �j@        G       H                    Z@*
;&���?             G@        ������������������������       �                      @        I       X                   po@�Ra����?             F@       J       U                   �_@�>4և��?             <@       K       T                    _@����X�?             ,@       L       S                    �?�θ�?
             *@       M       R                   0d@�q�q�?             "@       N       Q                   0c@      �?             @       O       P                    n@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        V       W                     M@@4և���?
             ,@       ������������������������       �        	             *@        ������������������������       �                     �?        ������������������������       �                     0@        Z       a                    �?�)�"*�?n             e@        [       `                   �d@$�q-�?             :@        \       _                   �n@r�q��?             (@        ]       ^                    c@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �        `            �a@        c       f                    �?�	j*D�?             *@        d       e                   �t@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        g       j                   �u@�����H�?             "@        h       i                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        l       w                    �?��T���?1            @R@       m       r       
             �?��-�=��?            �C@       n       q                    �F@��?^�k�?            �A@        o       p                    �D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @@        s       t                    @I@      �?             @        ������������������������       �                      @        u       v                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        x       y                    �?�!���?             A@        ������������������������       �                     (@        z       �                    b@      �?             6@       {       |                   �d@ҳ�wY;�?             1@        ������������������������       �                     @        }       �                   d@��
ц��?
             *@       ~       �       
             �?�z�G��?             $@              �       	          `ff�?      �?              @        �       �                   p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   i@ȵHPS!�?�            �s@        �       �       
             �?����˵�?F            �]@       �       �                    �?p�C��?7            �V@       ������������������������       �        +             R@        �       �                   @e@�KM�]�?             3@       �       �       
             �?�X�<ݺ?             2@        �       �                    �G@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     �?        �       �       	          033�?PN��T'�?             ;@       �       �                   @b@�}�+r��?
             3@       ������������������������       �                     *@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?B�1V���?            @h@        �       �                   �b@�s��:��?             C@       �       �                   `@���N8�?             5@       �       �                   @Z@�eP*L��?	             &@        ������������������������       �                     @        �       �                   �k@����X�?             @        ������������������������       �                     �?        �       �                   @`@r�q��?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?�t����?
             1@       �       �                    `@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?�8��8��?h            �c@        �       �                    �?r�q��?             B@        �       �                    �O@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �Z@�q�q�?             8@        ������������������������       �                     �?        �       �                    �?�㙢�c�?             7@       �       �                    �?�IєX�?             1@       ������������������������       �                     ,@        �       �                    @K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   @_@      �?             @        ������������������������       �                     �?        �       �                   �q@���Q��?             @        ������������������������       �                      @        �       �                     N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @i@�S���?M             ^@        ������������������������       �                      @        �       �                   �a@Xc!J�ƴ?L            �]@       �       �                   �c@��K2��?;            �W@       ������������������������       �        1            �S@        �       �                    �?��S�ۿ?
             .@       ������������������������       �                     (@        �       �                   r@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       	          033�?r�q��?             8@        ������������������������       �                     &@        �       �                   �b@�	j*D�?             *@        �       �                   �^@      �?             @        ������������������������       �                      @        �       �                    �K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?؇���X�?             @       ������������������������       �                     @        �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�Bp  ���>��?�,@��"�?��^Fb�?�׺Bs;�?G+�	�a�?r����<�?��y��y�?�a�a�?Cy�5��?^Cy�5�?UUUUUU�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?        �������?�������?              �?      �?                      �?Y�B��?��Moz��?�q�q�?��8��8�?              �?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�}�?��F���?�0���M�?�g *��?Q^Cy��?^Cy�5�?n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?""""""�?�������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?{	�%���?	�%����?]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?              �?      �?      �?                      �?      �?      �?              �?�������?�������?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?                      �?�b:��,�?�YLg1�?D��=��?��V!�n�?���,d!�?8��Moz�?              �?]t�E]�?]t�E�?�$I�$I�?�m۶m��?�m۶m��?�$I�$I�?ى�؉��?�؉�؉�?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?              �?      �?              �?                      �?n۶m۶�?�$I�$I�?      �?                      �?      �?        5���?ݾ�z�<�?�؉�؉�?;�;��?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        vb'vb'�?;�;��?      �?      �?              �?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �z��ի�?�B�
*�?�A�A�?}˷|˷�?�A�A�?_�_��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?�������?�������?      �?              �?      �?�������?�������?              �?�؉�؉�?�;�;�?333333�?ffffff�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?              �?        �؉�؉�?��N��N�?��/���?W'u_�?h�h��?��K��K�?              �?(�����?�k(���?�q�q�?��8��8�?�������?�������?      �?                      �?              �?      �?        h/�����?&���^B�?(�����?�5��P�?              �?UUUUUU�?�������?              �?      �?              �?      �?      �?                      �?��4l7��?���$2�?�k(���?��k(��?��y��y�?�a�a�?]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?�������?�������?�������?�������?              �?      �?              �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?        d!Y�B�?�7��Mo�?�?�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�����ݭ?""""""�?      �?        �pR�履?�؊���?W�+�Ʌ?��Q�٨�?              �?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?;�;��?vb'vb'�?      �?      �?      �?              �?      �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�-#hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKㅔh��B�8         b       	          ����?P��]��?�           ��@              +                    �?���a
�?�            �v@               
       
             �?��C���?[            �a@                     	          833�?R���Q�?3             T@       ������������������������       �        '            �O@               	                   �c@�t����?             1@                                  b@z�G�z�?             .@       ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                      @                                  @f@��6}��?(            �N@                                   �?     ��?             0@                     	          ����?�<ݚ�?             "@                                  Pb@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                   �H@����X�?             @                                  �^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               "                   �q@���V��?            �F@              !                   `p@�KM�]�?             C@                                 d@\-��p�?             =@                                  �K@�nkK�?             7@       ������������������������       �                     4@                                  �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                   �_@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        #       *                   �t@և���X�?             @       $       %                    �?      �?             @        ������������������������       �                     �?        &       '                     H@�q�q�?             @        ������������������������       �                     �?        (       )                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ,       M       
             �?>4և���?�             l@        -       <                   �a@b�2�tk�?%             K@       .       ;                    �? �Cc}�?             <@       /       :                    �?@�0�!��?             1@       0       1                    �?�θ�?	             *@        ������������������������       �                     �?        2       9                   p`@r�q��?             (@       3       8                   �b@�q�q�?             @       4       5                    @K@z�G�z�?             @        ������������������������       �                      @        6       7                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        =       H                   �e@�	j*D�?             :@       >       G                    �?��s����?             5@       ?       @                    �?�X�<ݺ?             2@        ������������������������       �                     @        A       B                   Pl@�8��8��?             (@        ������������������������       �                     @        C       D                    �H@r�q��?             @        ������������������������       �                     @        E       F       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        I       L                    �?z�G�z�?             @        J       K                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        N       _                   �t@�IєX�?g            @e@       O       X                    �?F|/ߨ�?d            @d@        P       S                    �?؇���X�?             5@       Q       R                   `b@�����H�?             2@       ������������������������       �                     0@        ������������������������       �                      @        T       W                    �?�q�q�?             @       U       V                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z       	            �?�k.s�׌?U            �a@       ������������������������       �        N             `@        [       ^                   p`@$�q-�?             *@        \       ]       	          pff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        `       a                   @c@      �?              @       ������������������������       �                      @        ������������������������       �                     @        c       �                   �c@������?�            w@       d       �                   Pr@���G�?�            t@       e       t                    �?lGts��?�            0q@        f       s       
             �?X�Cc�?             <@       g       n                   �^@��<b���?             7@        h       i                   �[@���Q��?             $@        ������������������������       �                     @        j       m                    �?z�G�z�?             @        k       l                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       p       	          ����?$�q-�?             *@       ������������������������       �                     "@        q       r                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        u       �                   P`@أ����?�            �n@        v       }                   �X@�t����?B            �]@        w       |                   pl@�	j*D�?             *@        x       {                    �?�q�q�?             @       y       z       	          `ff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ~       �                    a@0��_��?;            �Z@              �                    �?p��@���?/            @U@       �       �                    �?���C��?            �J@       �       �                    �K@@-�_ .�?            �B@       ������������������������       �                     ;@        �       �                    �L@z�G�z�?             $@        �       �                    ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?      �?	             0@        �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �       	             @�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @@        �       �                    @G@��s����?             5@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          `ff�?�����H�?
             2@        ������������������������       �                     "@        �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                   @_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   Pe@     �?S             `@        ������������������������       �                     E@        �       �                   �b@Du9iH��?9            �U@       �       �                    �?���J��?%            �I@       �       �                   �p@Pa�	�?            �@@       ������������������������       �                     ;@        �       �                    �L@r�q��?             @        ������������������������       �                     @        �       �                    �M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        �       �                   �e@؇���X�?            �A@        ������������������������       �                      @        �       �                    @�C��2(�?            �@@       �       �       
             �?      �?             @@       �       �       	          ����?(;L]n�?             >@        �       �                   �m@ףp=
�?             $@        ������������������������       �                     @        �       �                   �o@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          `ff�?8����?             G@        �       �                   �w@j���� �?             1@       �       �                    a@�θ�?
             *@       �       �                   �t@և���X�?             @       �       �                   @_@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?\-��p�?             =@        �       �       	          ���@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?�8��8��?             8@       ������������������������       �                     3@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?r�q��?             H@        �       �                   `T@d}h���?             ,@        ������������������������       �                      @        �       �                   d@�8��8��?             (@        �       �                   @`@z�G�z�?             @        ������������������������       �                     �?        �       �       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @b@�!���?             A@       �       �                    @�������?             >@       �       �                   �f@�q�q�?             5@       �       �       
             �?�<ݚ�?             2@        ������������������������       �                     @        �       �       	             @����X�?
             ,@       �       �                    @L@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  �h6n���?���� ��?�M5���?Ld���D�?g���Q��?L� &W�?333333�?333333�?              �?�������?�������?�������?�������?      �?                      �?              �?�!XG��?;ڼOq��?      �?      �?�q�q�?9��8���?      �?      �?      �?                      �?              �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        [�[��?�>�>��?�k(���?(�����?a����?�{a���?�Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        �m۶m��?%I�$I��?9��8���?�8��8��?۶m۶m�?%I�$I��?�������?ZZZZZZ�?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?              �?vb'vb'�?;�;��?z��y���?�a�a�?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?      �?              �?      �?                      �?�?�?�Hx�5�?�����H�?۶m۶m�?�$I�$I�?�q�q�?�q�q�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        "����?t�n��}?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?�On���?G:l��F�?�$RY���?�v����?�־a�?�<%�S��?�m۶m��?%I�$I��?��Moz��?��,d!�?�������?333333�?              �?�������?�������?      �?      �?              �?      �?              �?        ;�;��?�؉�؉�?              �?      �?      �?              �?      �?              �?        �KA���?���h�?�?<<<<<<�?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�V�9�&�?"5�x+��?�?�������?"5�x+��?\�琚`�?к����?S�n0E�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?      �?                      �?�q�q�?�q�q�?              �?      �?                      �?�a�a�?z��y���?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?     ��?              �?w�qGܱ?qG�w��?�?______�?|���?|���?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?        F]t�E�?]t�E�?      �?      �?�?�������?�������?�������?              �?      �?      �?      �?                      �?              �?      �?      �?              �?      �?              �?        8��Moz�?d!Y�B�?�������?ZZZZZZ�?ى�؉��?�؉�؉�?�$I�$I�?۶m۶m�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?                      �?�{a���?a����?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?              �?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?              �?        �������?�������?�������?�������?UUUUUU�?UUUUUU�?�q�q�?9��8���?              �?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ5�;5hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKͅ�h��B@3         ~       
             �?<���m�?�           ��@              Y                   �b@P@㞲��?           {@                                 �g@,sI�v�?�            �v@                                   �? ��+,��?Q            @_@                                   �?�:�]��?!            �I@       ������������������������       �                    �B@                                  Pa@����X�?
             ,@                                  �?X�<ݚ�?             "@       	       
                   0a@z�G�z�?             @        ������������������������       �                     @                                  �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        0            �R@               .                    �?t/*�?�            `m@                                   �?ҳ�wY;�?+             Q@                                  �[@b�2�tk�?             2@        ������������������������       �                     @                                   �?������?             .@                                  �N@      �?              @                                  @G@�q�q�?             @        ������������������������       �                     �?                                  Pb@z�G�z�?             @       ������������������������       �                     @                                  @q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                #                    @F@�-���?             I@        !       "                     D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        $       %                     L@�������?             F@        ������������������������       �                     .@        &       -       	             �?8^s]e�?             =@       '       ,                   �b@��.k���?             1@       (       )       	          ����?X�Cc�?	             ,@        ������������������������       �                     @        *       +                   @e@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             (@        /       :                   �[@�S-�?m            �d@        0       9                    �?D�n�3�?             3@       1       2       	             �?     ��?
             0@        ������������������������       �                     @        3       4                    �?�eP*L��?             &@        ������������������������       �                      @        5       8       	             �?�q�q�?             "@        6       7                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ;       J                   `\@@-�_ .�?a            �b@        <       E       	          ����?0��_��?#            �J@        =       @                   pm@���y4F�?             3@        >       ?                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        A       D                    �I@@4և���?             ,@        B       C                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        F       G                    �?г�wY;�?             A@       ������������������������       �                     =@        H       I                    �Q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        K       P                    �?�==Q�P�?>            �W@       L       M                    f@��'�`�?6            �T@       ������������������������       �        2            �S@        N       O                   �s@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        Q       X                   �s@r�q��?             (@       R       S                   �`@�C��2(�?             &@       ������������������������       �                     @        T       U                    n@z�G�z�?             @        ������������������������       �                      @        V       W                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        Z       g                    �?b1<+�C�?/            @R@        [       `                   �^@���@��?            �B@        \       _                    �?      �?             ,@       ]       ^       	          ����?�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        a       f                    �?�nkK�?             7@        b       e                   �c@�8��8��?             (@        c       d                    b@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        h       w       	          033�?X�<ݚ�?             B@       i       j                    @H@�	j*D�?             :@        ������������������������       �                     $@        k       l       
             �?      �?             0@        ������������������������       �                      @        m       n                   �h@և���X�?
             ,@        ������������������������       �                     @        o       p                   �l@�eP*L��?             &@        ������������������������       �                     @        q       t                    a@      �?              @        r       s                   e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        u       v                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        x       }                    �N@z�G�z�?             $@       y       |                    �?�����H�?             "@       z       {                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               �       	          ����?D� r�?�            �r@       �       �                    �?�K�w���?�            `l@        �       �                   �b@6��f�?.            @S@       �       �                    �?���7�?             F@       �       �       	            �?�(\����?             D@       ������������������������       �                     A@        �       �                    V@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �Z@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �i@4���C�?            �@@        �       �                   �e@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�	j*D�?             :@       �       �                    �?���N8�?             5@       �       �                   �q@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �l@ףp=
�?             $@        ������������������������       �                     @        �       �       	          ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �l@���Q��?             @        ������������������������       �                     �?        �       �                     M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	            �?�}��L�?g            �b@       �       �                   0a@ ��U��?c            �a@       ������������������������       �        I            @Z@        �       �                   �c@�?�|�?            �B@       �       �                   �a@�IєX�?             1@        �       �                   @c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             &@        ������������������������       �                     4@        �       �                    �M@      �?              @        �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?,            �R@       �       �                   @b@�I�w�"�?             C@       �       �                   ht@HP�s��?             9@       �       �                    �H@ �q�q�?             8@        �       �                   �Z@r�q��?             @        ������������������������       �                     @        �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                     �?        �       �       	             �?��
ц��?             *@       �       �                   �s@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    ]@�<ݚ�?             B@        ������������������������       �                     @        �       �                    �?6YE�t�?            �@@        ������������������������       �                     ,@        �       �                    �?�d�����?             3@        ������������������������       �                      @        �       �                    �?@�0�!��?             1@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       	             @؇���X�?             ,@       �       �                    j@$�q-�?             *@       �       �                   0i@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ���>��?�,@��"�?t�>v�H�?#Up�ѭ�?��I��I�?l�l��?����Mb�?`��"���?�?}}}}}}�?              �?�$I�$I�?�m۶m��?�q�q�?r�q��?�������?�������?      �?              �?      �?              �?      �?                      �?              �?              �?W�+���?�;����?�������?�������?�8��8��?9��8���?              �?wwwwww�?�?      �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?      �?                      �?              �?      �?        �p=
ף�?�G�z��?UUUUUU�?UUUUUU�?              �?      �?        /�袋.�?t�E]t�?              �?	�=����?|a���?�������?�?%I�$I��?�m۶m��?              �?/�袋.�?F]t�E�?      �?                      �?              �?              �?J���冸?���A#��?(������?l(�����?      �?      �?              �?]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        к����?S�n0E�?�V�9�&�?"5�x+��?(������?6��P^C�?333333�?�������?      �?                      �?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?�?�?              �?�������?�������?              �?      �?        �a�+�?��%N��?��k���?1P�M��?              �?�������?�������?              �?      �?        UUUUUU�?�������?F]t�E�?]t�E�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        Ĉ#F��?�;w�ܹ�?к����?L�Ϻ��?      �?      �?ffffff�?333333�?              �?      �?                      �?d!Y�B�?�Mozӛ�?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?                      �?              �?              �?r�q��?�q�q�?vb'vb'�?;�;��?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?              �?t�E]t�?]t�E�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?�������?�������?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        ���w'�?٥Q �c�?�hAjv�?����L�?g�'�Y�?�cj`��?�.�袋�?F]t�E�?333333�?�������?      �?        �������?UUUUUU�?              �?      �?              �?      �?              �?      �?        m��&�l�?'�l��&�?�$I�$I�?۶m۶m�?              �?      �?        vb'vb'�?;�;��?�a�a�?��y��y�?]t�E]�?F]t�E�?      �?                      �?�������?�������?      �?              �?      �?      �?                      �?�������?333333�?      �?              �?      �?              �?      �?        �_,�Œ�?O贁N�?���RO��?��V�|?      �?        *�Y7�"�?к����?�?�?�������?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?      �?              �?      �?              �?              �?      �?�5��P�?����k�?{�G�z�?q=
ףp�?UUUUUU�?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �;�;�?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?              �?        9��8���?�q�q�?              �?'�l��&�?e�M6�d�?      �?        Cy�5��?y�5���?              �?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?�������?�������?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJi4�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK煔h��B�9         v       	          033�?��;/M�?�           ��@              E                    �?r�q��?�             x@               4                    @M@�C���?f            �d@                                  �?r�q��?H             ^@                     
             �?.�W����?0            �R@                                   �?H%u��?             9@                                 �_@؇���X�?             5@       ������������������������       �        	             .@        	       
       	          @33�?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                   Z@HP�s��?              I@        ������������������������       �                      @                                   �? �q�q�?             H@        ������������������������       �                     "@                                  �_@�7��?            �C@                                  `\@؇���X�?             @       ������������������������       �                     @                                  �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                      	          ����?      �?             @@       ������������������������       �                     ?@        ������������������������       �                     �?               /                    �?�L�lRT�?            �F@                                 Pg@4���C�?            �@@        ������������������������       �                     @               $                    ^@��
ц��?             :@               #                   �[@�<ݚ�?             "@                                  `k@      �?             @        ������������������������       �                     �?        !       "                    @L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        %       (                   @`@�t����?	             1@        &       '                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        )       .       
             �?r�q��?             (@       *       +       	          ����?      �?             @        ������������������������       �                     �?        ,       -                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        0       3                    b@r�q��?             (@       1       2                   Xp@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        5       D                   `f@�㙢�c�?             G@       6       A       	          833�?���V��?            �F@       7       8       
             �?     ��?             @@       ������������������������       �                     4@        9       @                    `Q@      �?             (@       :       ?                    �N@      �?              @       ;       >                   �b@����X�?             @       <       =                   �e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        B       C                   @]@�	j*D�?             *@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     �?        F       g                    �?Rԅ5l�?�            @k@       G       L                    �?�LQ�1	�?             g@        H       I                   r@`׀�:M�?1            �R@       ������������������������       �        )             P@        J       K       
             �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        M       X       
             �?p��*�?N            �[@        N       U                    �?�X����?             6@        O       T                     N@�q�q�?             "@       P       Q       
             �?؇���X�?             @        ������������������������       �                      @        R       S                     C@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        V       W                    �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �        
             (@        Y       b       	            �?�C��2(�?=             V@       Z       _                    �N@ �\���?6            �S@       [       \                    @L@P�Lt�<�?4             S@       ������������������������       �        0            �P@        ]       ^                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        `       a                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        c       f                   a@X�<ݚ�?             "@       d       e                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        h       q       
             �?j���� �?             A@        i       j       	          ����?     ��?	             0@       ������������������������       �                     "@        k       l                    �H@և���X�?             @        ������������������������       �                      @        m       n                   `_@z�G�z�?             @        ������������������������       �                      @        o       p                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        r       u                    �?�X�<ݺ?             2@        s       t                   �`@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        w       �                    �?���lv	�?�            �u@        x       �                   �a@��o	��?)             M@       y       �                   `a@�D����?             E@       z       �                    �?П[;U��?             =@       {       |       
             �?�q�q�?             2@        ������������������������       �                      @        }       �                    �?      �?
             0@       ~                            N@$�q-�?             *@       ������������������������       �                     $@        �       �                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�C��2(�?
             &@       ������������������������       �        	             $@        ������������������������       �                     �?        �       �                   �a@$�q-�?	             *@       ������������������������       �                     &@        �       �       	          033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?      �?             0@       ������������������������       �        
             ,@        ������������������������       �                      @        �       �                    �F@�)�0���?�            @r@        �       �                    �?�q�q�?             8@        �       �                    �?�q�q�?             "@       �       �       	             @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �_@�r����?
             .@        ������������������������       �                      @        �       �                    b@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �z@,T\��?�            �p@       �       �                    �?���C��?�            �p@       �       �       	          ����?�8��8��?�             k@        �       �                    �?�:pΈ��?<             Y@        �       �                   pr@�I�w�"�?             C@       �       �       
             �?tk~X��?             B@        �       �                   �^@      �?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �       	             �?$�q-�?             :@        �       �                    �?      �?              @        �       �                   �q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                      @        �       �                   P`@6uH���?)             O@        �       �                   �X@r�q��?             8@        �       �                    �K@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    ]@�X�<ݺ?             2@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                    @N@�q�q�?             @       �       �                    Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             (@        �       �                   P`@P�Lt�<�?             C@       ������������������������       �                     =@        �       �       
             �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                     R@XB���?H             ]@       �       �                    c@ T���v�?F            @\@       �       �                   �c@@3����?B             [@       �       �                    \@�L��ȕ?8            @W@        �       �                   �_@ ���J��?            �C@        �       �                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �        $             K@        �       �                    �?��S�ۿ?
             .@        �       �                   p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                   pc@z�G�z�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `b@ \� ���?!            �H@       �       �                   ``@R���Q�?             D@       �       �                    `@      �?             8@       �       �                    @P@�KM�]�?             3@       ������������������������       �                     .@        �       �                   �]@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     0@        �       �                   0a@�q�q�?             "@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  �X�5��?�S�$e�?UUUUU�?UUUUU��?�!�%�?	o4u~��?UUUUUU�?UUUUUU�?贁N��?0��b�/�?���Q��?)\���(�?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?q=
ףp�?{�G�z�?              �?�������?UUUUUU�?      �?        ��[��[�?�A�A�?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?      �?      �?                      �?l�l��?�I��I��?'�l��&�?m��&�l�?              �?�;�;�?�؉�؉�?�q�q�?9��8���?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?�������?333333�?      �?                      �?�������?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?�$I�$I�?�m۶m��?              �?      �?                      �?d!Y�B�?�7��Mo�?�>�>��?[�[��?      �?      �?              �?      �?      �?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?              �?              �?                      �?;�;��?vb'vb'�?              �?      �?              �?        ���d	l�?�d	l�O�?��Moz��?Y�B��?��L��?к����?      �?        �������?�������?              �?      �?        O	� O�?��7�}��?]t�E]�?�E]t��?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?                      �?;�;��?�؉�؉�?      �?                      �?]t�E�?F]t�E�?���7a�?�3���?���k(�?(�����?      �?        9��8���?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        r�q��?�q�q�?�������?�������?              �?      �?              �?        �������?ZZZZZZ�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ��8��8�?�q�q�?�������?�������?      �?                      �?      �?        L�w�Z��?�bSi��?������?���{�?�0�0�?z��y���?��=���?�{a���?UUUUUU�?UUUUUU�?              �?      �?      �?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?]t�E�?              �?      �?        �؉�؉�?;�;��?      �?              �?      �?              �?      �?              �?      �?              �?      �?        �?~���?8p����?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?              �?�?�������?              �?�$I�$I�?�m۶m��?              �?      �?        "=P9���?\�՘H�?"5�x+��?\�琚`�?UUUUUU�?UUUUUU�?�Q����?��Q���?�5��P�?����k�?9��8���?r�q��?      �?      �?              �?      �?        ;�;��?�؉�؉�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        ��RJ)��?k���Zk�?UUUUUU�?�������?      �?      �?              �?      �?        �q�q�?��8��8�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?(�����?���k(�?              �?�q�q�?�q�q�?              �?      �?        �{a���?GX�i���?4��A�/�?6h�e�&�?h/�����?���Kh�?X`��?��~���?�A�A�?��-��-�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�?�������?      �?      �?      �?                      �?              �?�������?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        և���X�?
^N��)�?333333�?333333�?      �?      �?(�����?�k(���?              �?      �?      �?      �?                      �?�������?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ThG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKŅ�h��B@1         �       
             �?� 07��?�           ��@              e                   �b@�}
��?	           z@              <                   �`@��<���?�            �u@                                  �c@�����?b            `b@               
                   �X@��Y��]�?            �D@               	       	             �?z�G�z�?             @                                  @M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     B@               7       	          `ff�?r�0p�?D            �Z@              "                    �?���|���?/            @S@                      	          @33�?h+�v:�?             A@                                   �?�<ݚ�?             "@       ������������������������       �                     @                                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  @l@�+e�X�?             9@        ������������������������       �                     @                                   �K@�q�q�?             2@        ������������������������       �                      @                                  �T@���Q��?             $@        ������������������������       �                      @               !                   �b@      �?              @                                  �o@���Q��?             @                                 �\@�q�q�?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        #       .                    �?�T|n�q�?            �E@       $       %                   0i@�C��2(�?            �@@        ������������������������       �                     �?        &       -                    @      �?             @@       '       (                   @_@�g�y��?             ?@       ������������������������       �                     6@        )       ,                    `@�����H�?             "@        *       +                    Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        /       0                    �?���Q��?             $@        ������������������������       �                     @        1       6                   �l@և���X�?             @       2       5                   �j@���Q��?             @       3       4       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        8       ;                    �J@XB���?             =@        9       :                    @J@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        =       d                    �R@������?x            �h@       >       S                    �? ���v��?w            �h@       ?       P                    `R@      �?_             d@       @       O                    �? ���J��?\            �c@       A       H                   �h@�94�s0�?D            �\@        B       G                   Pb@HP�s��?             9@       C       D                   �_@ �q�q�?             8@       ������������������������       �                     3@        E       F                    �I@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        I       J                    @K@����?�?4            �V@        ������������������������       �                     C@        K       N       	          ����? ��WV�?             J@        L       M                     M@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     H@        ������������������������       �                    �D@        Q       R                   �p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        T       a                    �Q@�?�'�@�?             C@       U       \                   �e@�C��2(�?            �@@       V       W                   a@ ��WV�?             :@       ������������������������       �                     3@        X       Y                    �?؇���X�?             @       ������������������������       �                     @        Z       [                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ]       ^                    �?����X�?             @        ������������������������       �                     @        _       `                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        b       c                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        f       g                    @C@`��_��?/            �Q@        ������������������������       �                      @        h       i                    @G@X�<ݚ�?*            �O@        ������������������������       �        
             ,@        j       o                    @H@և���X�?             �H@        k       n       	          hff�?؇���X�?             ,@        l       m       	          ����?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        p       s                    �J@�xGZ���?            �A@        q       r                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        t       u                   0c@X�<ݚ�?             ;@        ������������������������       �                     @        v       }                   d@      �?             8@       w       x                    �?z�G�z�?             .@        ������������������������       �                     @        y       z                    @M@�z�G��?             $@       ������������������������       �                     @        {       |                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ~       �                    �?�q�q�?             "@              �                     L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   `R@ ���:�?�            �s@        �       �                     E@X�<ݚ�?             ;@        ������������������������       �                     @        �       �       	          hff�?      �?             8@        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          `ff�?@�0�!��?             1@       �       �                   `b@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                    �?���Q��?             @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?��ϭ�*�?�             r@       �       �                    @L@؝�x�O�?�            �p@       �       �                    �?��6�.ӯ?~            @k@        �       �                    �H@r�q��?             >@       �       �                   @^@�t����?             1@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     *@        �       �                    �?��K2��?k            �g@        �       �       	          433�?�X�<ݺ?             B@       �       �                   �l@�g�y��?             ?@        ������������������������       �        	             .@        �       �                   0c@      �?
             0@       ������������������������       �                     *@        �       �                   0d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?z�G�z�?             @        �       �                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        S             c@        �       �       	          033@��x_F-�?!            �I@       �       �       	          ����?��E�B��?            �G@       �       �                   d@`2U0*��?             9@       ������������������������       �                     ,@        �       �                   `c@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �?�GN�z�?             6@        ������������������������       �                     @        �       �                    �M@�t����?
             1@        �       �                    e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        �       �                   �r@�ՙ/�?             5@       �       �                    �?������?             1@       �       �       	          ����?X�<ݚ�?             "@       �       �                   �b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�b���      h�h)h,K ��h.��R�(KK�KK��hb�BP  ������?
��,@��?��T�?��;?�*�?Z/`��U�?���E5�?����X�?^N��)x�?������?8��18�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?oe�Cj��?HM0��>�?F]t�E�?]t�E]�?�������?xxxxxx�?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?        R���Q�?���Q��?      �?        UUUUUU�?UUUUUU�?      �?        �������?333333�?      �?              �?      �?�������?333333�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?              �?6eMYS��?���)k��?F]t�E�?]t�E�?      �?              �?      �?�B!��?��{���?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?333333�?              �?�$I�$I�?۶m۶m�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �{a���?GX�i���?      �?      �?              �?      �?                      �?���/M�?�n-;�?1ogH�۩?�y;Cb�?      �?      �?�A�A�?��-��-�?���ϡ?��%���?{�G�z�?q=
ףp�?UUUUUU�?�������?              �?�������?�������?      �?                      �?      �?        l�l��?��I��I�?              �?;�;��?O��N���?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?        y�5���?������?F]t�E�?]t�E�?;�;��?O��N���?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?�������?333333�?      �?                      �?      �?        ��ۥ���?6��9�?              �?r�q��?�q�q�?      �?        ۶m۶m�?�$I�$I�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?�_�_�?�A�A�?      �?      �?      �?                      �?�q�q�?r�q��?      �?              �?      �?�������?�������?              �?333333�?ffffff�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �7W$O��?!�n�&�?�q�q�?r�q��?      �?              �?      �?۶m۶m�?�$I�$I�?      �?                      �?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?      �?      �?      �?                      �?              �?����=�?|a���?�� ;J��?�b�'�-�?���A���?��p�?�������?UUUUUU�?�������?�������?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?              �?        ��Q�٨�?W�+�Ʌ?��8��8�?�q�q�?��{���?�B!��?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?              �?      �?              �?              �?        �������?�?�l�w6��?AL� &W�?���Q��?{�G�z�?      �?        ]t�E�?F]t�E�?      �?                      �?�袋.��?]t�E�?      �?        �������?�������?UUUUUU�?�������?              �?      �?              �?                      �?�<��<��?�a�a�?xxxxxx�?�?r�q��?�q�q�?�������?UUUUUU�?      �?                      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ5�R/hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@>         �       
             �?T8���?�           ��@              S                    �?Z�K��?            z@                                  �F@������?�            �q@               	                    Z@      �?             <@                      	             @�q�q�?             @                                 �o@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        
              	          ����?��2(&�?             6@        ������������������������       �                     $@                                  �a@      �?             (@                     	          ����?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @               F       	          pff�?�L���?�            0p@              C                   �u@T����?g            @c@              B                    �?,I�e���?e            �b@                                 `\@�ջ����?G             Z@                                   �K@X�<ݚ�?             "@                                  �k@      �?             @        ������������������������       �                      @                                   �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �M@z�G�z�?             @        ������������������������       �                     @                      	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                '                    @K@�j�@�?@            �W@        !       "                    @J@P�Lt�<�?             C@       ������������������������       �                     9@        #       &                    �?$�q-�?             *@        $       %       	          hff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        (       ;                   pb@F�t�K��?$            �L@       )       *       	          ����?8�Z$���?              J@        ������������������������       �                     .@        +       0                    �?���@��?            �B@        ,       -       
             �?�q�q�?             @        ������������������������       �                      @        .       /       	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        1       2       	          hff�?��� ��?             ?@        ������������������������       �                     �?        3       6       	          ����?ףp=
�?             >@        4       5                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        7       8                    �?�>����?             ;@       ������������������������       �        	             4@        9       :                   ``@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        <       =                   0a@���Q��?             @        ������������������������       �                      @        >       ?                    �?�q�q�?             @        ������������������������       �                     �?        @       A                    @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �G@        D       E                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        G       R                   �a@P�c0"�?D            @Z@       H       I                   8p@0�,���?+            �P@       ������������������������       �                    �H@        J       O                   pa@�����H�?             2@       K       N                   �_@@4և���?             ,@       L       M                   �^@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        P       Q                   `a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     C@        T       �       	          `ff�?��>^�?Q             `@       U       n                   �a@և���X�?@            �X@        V       a       	          ����?��x_F-�?             �I@       W       X                    �?��a�n`�?             ?@        ������������������������       �                     �?        Y       `                    �?��S�ۿ?             >@       Z       _                    j@�����H�?	             2@       [       \                   @`@����X�?             @       ������������������������       �                     @        ]       ^                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     (@        b       m                   �`@��Q��?             4@       c       j       	          ����?������?             1@       d       i       	             �?      �?              @       e       h                   �]@����X�?             @       f       g                    @Q@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        k       l                    �Q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        o       r                   `h@(���@��?             �G@        p       q       	          033�?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        s       �                    �P@���?            �D@       t       �                    @K@>A�F<�?             C@       u       �                    �?����X�?             5@       v       w                   pk@@�0�!��?             1@        ������������������������       �                     @        x       y                    �?�z�G��?
             $@        ������������������������       �                     @        z       �                   �e@և���X�?             @       {       |                   �\@���Q��?             @        ������������������������       �                     �?        }       ~                   0c@      �?             @        ������������������������       �                     �?               �                   pd@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �l@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   a@�IєX�?	             1@       ������������������������       �                     "@        �       �                    @      �?              @        ������������������������       �                     @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��� ��?             ?@       �       �                    �F@�<ݚ�?
             2@        ������������������������       �                      @        �       �                    �?      �?	             0@        ������������������������       �                     �?        �       �                    �?��S�ۿ?             .@       ������������������������       �                     *@        �       �                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    �?�� �?�            �s@       �       �                    @L@d/�@7�?�             q@       �       �                    �?88��M�?�            �j@        �       �                   @\@�>4և��?             <@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@�8��8��?             8@        �       �                    @H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             2@        �       �       	          ����?Hn�.P��?o            @g@       �       �                   @E@@�?�c�?b            �d@        �       �                    �B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��z*�o�?^            �c@       �       �                    ]@     ��?M             `@        �       �                   �c@���}<S�?             7@       ������������������������       �                     .@        �       �                    �?      �?              @       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        >            @Z@        ������������������������       �                     ?@        �       �                    �?���!pc�?             6@        �       �                   `T@�q�q�?             "@        ������������������������       �                     @        �       �                   pe@���Q��?             @       �       �                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        �       �                   �a@d��0u��?$             N@        �       �       	          (33�?"pc�
�?             6@       �       �                   @\@�IєX�?             1@        �       �       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�\��N��?             C@        �       �                   �_@X�Cc�?             ,@        ������������������������       �                     @        �       �                     O@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �L@r�q��?             8@        ������������������������       �                     @        �       �                   Pb@D�n�3�?             3@        ������������������������       �                     @        �       �                    �?     ��?             0@        �       �                   `c@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ��� @r�q��?             (@       �       �                   ps@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     M@8�A�0��?             F@       �       �                    �?�q�q�?             8@        ������������������������       �                     @        �       �                   b@j���� �?             1@       �       �                    �F@      �?              @        ������������������������       �                     �?        �       �                   �Z@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �C@�����H�?             "@        ������������������������       �                     @        �       �                     G@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?             4@        ������������������������       �                     �?        �       �                   �]@�S����?             3@        �       �                    �?���Q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �^@@4և���?	             ,@        �       �                    �?      �?             @       �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  6n����?�� ���?O��N���?��N��N�?������?�|����?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        t�E]t�?��.���?              �?      �?      �?�������?�������?      �?                      �?      �?        L�Ϻ��?}���g�?qV~B���?25�wL�?�Hs�9Ҽ?�q˸e�?�N��N��?O��N���?r�q��?�q�q�?      �?      �?              �?      �?      �?      �?                      �?�������?�������?      �?              �?      �?              �?      �?        �a�+�?T��8��?(�����?���k(�?              �?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?              �?:��,���?1��t��?;�;��?;�;��?              �?к����?L�Ϻ��?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�B!��?�{����?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?h/�����?�Kh/��?              �?�$I�$I�?�m۶m��?      �?                      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        8�8��??�c?�c�?g��1��?Ez�rv�?              �?�q�q�?�q�q�?�$I�$I�?n۶m۶�?UUUUUU�?�������?              �?      �?                      �?      �?      �?              �?      �?                      �?�%mI[��?&mI[Җ�?۶m۶m�?�$I�$I�?�?�������?�c�1Ƹ?�s�9��?      �?        �?�������?�q�q�?�q�q�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?ffffff�?�������?�?xxxxxx�?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?              �?              �?        �q�q�?�q�q�?              �?      �?              �?        W�+���?R�٨�l�?UUUUUU�?�������?              �?      �?        28��1�?8��18�?������?Cy�5��?�m۶m��?�$I�$I�?ZZZZZZ�?�������?      �?        ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?�?�?      �?              �?      �?      �?              �?      �?      �?                      �?              �?�B!��?�{����?�q�q�?9��8���?      �?              �?      �?      �?        �?�������?              �?      �?      �?      �?                      �?              �?��N���?�{mĺ��?�ǭ��?��;�H��?+J�#��?����f��?�$I�$I�?�m۶m��?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        t�9�s�?�c�1ƨ?jW�v%j�?��+Q��?�������?�������?              �?      �?        |mĺ���?��N�?     ��?      �?ӛ���7�?d!Y�B�?      �?              �?      �?      �?              �?      �?              �?      �?              �?              �?        F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?              �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        DDDDDD�?wwwwww�?/�袋.�?F]t�E�?�?�?�������?�������?      �?                      �?      �?        �������?333333�?      �?                      �?y�5���?�5��P�?%I�$I��?�m۶m��?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?l(�����?(������?              �?      �?      �?      �?      �?      �?      �?      �?                      �?              �?�������?UUUUUU�?]t�E�?F]t�E�?      �?                      �?              �?/�袋.�?颋.���?�������?�������?      �?        ZZZZZZ�?�������?      �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?        �q�q�?�q�q�?              �?�������?�������?      �?                      �?�������?�������?      �?        ^Cy�5�?(������?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?n۶m۶�?      �?      �?      �?      �?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�%hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKم�h��B@6         �       
             �?.��X~��?�           ��@                                 �a@g\�i�?           0z@               
                    �?`Jj��?M             _@              	                    �Q@(;L]n�?7            �V@                                 `X@�x�E~�?6            @V@                                  �W@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �        .            �S@        ������������������������       �                     �?                                   �?��hJ,�?             A@       ������������������������       �                     8@                                  @_@      �?             $@        ������������������������       �                      @                      	          `ff�?      �?              @        ������������������������       �                      @                      	             @r�q��?             @        ������������������������       �                     @                                  c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               m       	          pff�?v���~�?�            pr@              R                   Pa@>�V�n��?|             g@              5                    �?V�s�s�?P            �^@               .                    �?�L�lRT�?            �F@                                  �?�n`���?             ?@        ������������������������       �                     @               #                    �?      �?             8@               "                    �?      �?              @                                 `m@�q�q�?             @        ������������������������       �                     �?                !       	          `ff�?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        $       %                   �]@      �?             0@        ������������������������       �                     @        &       '                   `X@z�G�z�?             $@        ������������������������       �                     �?        (       -                   �b@�����H�?             "@        )       ,                    @L@      �?             @       *       +       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        /       0                   �`@����X�?	             ,@       ������������������������       �                     @        1       2                    l@և���X�?             @        ������������������������       �                      @        3       4                   (p@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        6       E                    �?��cv�?3            @S@       7       8                     L@8��8���?!             H@       ������������������������       �                     ;@        9       D                   r@�q�q�?             5@       :       ;       
             �?�d�����?             3@        ������������������������       �                      @        <       A                    �?�t����?
             1@        =       >                    �M@և���X�?             @        ������������������������       �                     @        ?       @                   �\@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        B       C                    �L@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        F       I                   �a@�f7�z�?             =@        G       H                   �\@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        J       O                     I@�d�����?             3@        K       L                   `]@�q�q�?             @        ������������������������       �                     @        M       N                    l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        P       Q       	          ����?$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        S       d                    �?�<ݚ�?,            �O@       T       ]                   �a@��0{9�?!            �G@        U       \                    b@�q�q�?             .@       V       [                    �?r�q��?	             (@       W       Z       	             �?z�G�z�?             $@        X       Y                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ^       _                    �E@      �?             @@        ������������������������       �                     �?        `       a                   `f@�g�y��?             ?@       ������������������������       �                     =@        b       c                   �s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        e       l                    �?     ��?             0@       f       g                    �?��
ц��?	             *@        ������������������������       �                     @        h       i                    �N@      �?              @       ������������������������       �                     @        j       k                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        n       o                   �Z@X�;�^o�?G            �[@        ������������������������       �                      @        p       q                   �j@�����H�?F             [@        ������������������������       �                     4@        r                           �?��2(&�?9             V@        s       t                   �^@      �?             <@        ������������������������       �                     @        u       v                    _@�q�q�?             5@        ������������������������       �                      @        w       |                   Pn@�d�����?             3@        x       y                    �?�q�q�?             @        ������������������������       �                      @        z       {                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        }       ~                    �?$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �                    c@�8��8��?(             N@       �       �                   �c@ ,��-�?'            �M@       �       �                    �? �q�q�?!             H@        ������������������������       �                     �?        �       �       	          033@`Ql�R�?             �G@       ������������������������       �                     >@        �       �                   �_@�IєX�?             1@        �       �                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        �       �                   r@"pc�
�?             &@        ������������������������       �                     @        �       �       
             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @c@4�2%ޑ�?�            �s@        �       �                    �?���c�H�?            �H@       �       �       	          @33�?
j*D>�?             :@        �       �                   p`@z�G�z�?             $@       ������������������������       �                     @        �       �                   �]@���Q��?             @        ������������������������       �                      @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?     ��?             0@        ������������������������       �                     @        �       �                    �?�θ�?             *@        ������������������������       �                      @        �       �                    �I@���Q��?             @        ������������������������       �                     �?        �       �                    �M@      �?             @        ������������������������       �                     �?        �       �       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        �       �                    �?��F���?�            �p@        �       �                    s@Ћ����?:            �T@       ������������������������       �        ,             N@        �       �                    �?��2(&�?             6@        �       �                    �?�q�q�?             "@        ������������������������       �                      @        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        �       �       	          833�?lK���?r             g@       �       �                    @L@�W����?Z            �a@       �       �                    �?�T�~~4�?H            @]@        �       �                    �?�>����?             ;@       �       �                   �\@���}<S�?             7@        �       �                   �g@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     @        ������������������������       �        6            �V@        �       �                   0c@z�G�z�?             9@       �       �                   �_@�X�<ݺ?             2@        �       �                   �^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             .@        �       �                    �?և���X�?             @       �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?և���X�?             E@       �       �                    d@�X����?             6@       �       �                   ``@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �       	             �?�eP*L��?             &@        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                   ``@�q�q�?             @        ������������������������       �                      @        �       �                   �e@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?R���Q�?             4@       �       �                    �?z�G�z�?	             .@       ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��� ���?���o���?���mD0�?����3�?�B!��?���{��?�?�������?p�\��?����G�?F]t�E�?/�袋.�?              �?      �?                      �?      �?        �������?KKKKKK�?              �?      �?      �?              �?      �?      �?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �7@Z���?;��ҫ6�?�r�4�-�?�F��*i�?q�����?G��).�?�I��I��?l�l��?�9�s��?�c�1��?      �?              �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?              �?      �?      �?        �������?�������?              �?�q�q�?�q�q�?      �?      �?      �?      �?              �?      �?              �?              �?        �$I�$I�?�m۶m��?              �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?                      �?��O����?��;��?�������?UUUUUU�?              �?UUUUUU�?UUUUUU�?y�5���?Cy�5��?              �?�������?�������?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?        �������?�������?      �?                      �?      �?        O#,�4��?a���{�?333333�?ffffff�?      �?                      �?Cy�5��?y�5���?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?;�;��?      �?                      �?�q�q�?9��8���?L� &W�?m�w6�;�?UUUUUU�?UUUUUU�?UUUUUU�?�������?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?              �?      �?      �?        �B!��?��{���?              �?      �?      �?              �?      �?              �?      �?�;�;�?�؉�؉�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?J��yJ�?�־a��?      �?        �q�q�?�q�q�?              �?t�E]t�?��.���?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        y�5���?Cy�5��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ;�;��?�؉�؉�?              �?      �?        UUUUUU�?UUUUUU�?'u_[�?[4���?UUUUUU�?�������?      �?        W�+�ɕ?}g���Q�?              �?�?�?      �?      �?      �?                      �?              �?F]t�E�?/�袋.�?              �?�������?333333�?      �?                      �?      �?        �������?�A�A�?/�����?4և����?;�;��?b'vb'v�?�������?�������?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?�؉�؉�?ى�؉��?              �?333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?��9����?�d\�?ԮD�J��?��+Q��?      �?        ��.���?t�E]t�?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?        �Mozӛ�?Y�B���?�́D+l�?�'�K=�??�s?�s�?���?�Kh/��?h/�����?ӛ���7�?d!Y�B�?333333�?�������?              �?      �?              �?              �?              �?        �������?�������?��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?�E]t��?]t�E]�?]t�E�?F]t�E�?              �?      �?        ]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        333333�?333333�?�������?�������?              �?      �?                      �?�t�bubhhubehhub.